// DSCH 3.5
// 29-11-2022 15:26:02
// C:\Users\savit\Downloads\BoothMultiplier.sch

module BoothMultiplier( MC3,MC2,MC1,MC0,MP3,MP2,MP1,MP0,
 PROD7,PROD6,PROD5,PROD4,PROD3,PROD2,PROD1,PROD0);
 input MC3,MC2,MC1,MC0,MP3,MP2,MP1,MP0;
 output PROD7,PROD6,PROD5,PROD4,PROD3,PROD2,PROD1,PROD0;
 wire w18,w19,w20,w21,w22,w23,w24,w25;
 wire w26,w27,w28,w29,w30,w31,w32,w33;
 wire w34,w35,w36,w37,w38,w39,w40,w41;
 wire w42,w43,w44,w45,w46,w47,w48,w49;
 wire w50,w51,w52,w53,w54,w55,w56,w57;
 wire w58,w59,w60,w61,w62,w63,w64,w65;
 wire w66,w67,w68,w69,w70,w71,w72,w73;
 wire w74,w75,w76,w77,w78,w79,w80,w81;
 wire w82,w83,w84,w85,w86,w87,w88,w89;
 wire w90,w91,w92,w93,w94,w95,w96,w97;
 wire w98,w99,w100,w101,w102,w103,w104,w105;
 wire w106,w107,w108,w109,w110,w111,w112,w113;
 wire w114,w115,w116,w117,w118,w119,w120,w121;
 wire w122,w123,w124,w125,w126,w127,w128,w129;
 wire w130,w131,w132,w133,w134,w135,w136,w137;
 wire w138,w139,w140,w141,w142,w143,w144,w145;
 wire w146,w147,w148,w149,w150,w151,w152,w153;
 wire w154,w155,w156,w157,w158,w159,w160,w161;
 wire w162,w163,w164,w165,w166,w167,w168,w169;
 wire w170,w171,w172,w173,w174,w175,w176,w177;
 wire w178,w179,w180,w181,w182,w183,w184,w185;
 wire w186,w187,w188,w189,w190,w191,w192,w193;
 wire w194,w195,w196,w197,w198,w199,w200,w201;
 wire w202,w203,w204,w205,w206,w207,w208,w209;
 wire w210,w211,w212,w213,w214,w215,w216,w217;
 wire w218,w219,w220,w221,w222,w223,w224,w225;
 wire w226,w227,w228,w229,w230,w231,w232,w233;
 wire w234,w235,w236,w237,w238,w239,w240,w241;
 wire w242,w243,w244,w245,w246,w247,w248,w249;
 wire w250,w251,w252,w253,w254,w255,w256,w257;
 wire w258,w259,w260,w261,w262,w263,w264,w265;
 wire w266,w267,w268,w269,w270,w271,w272,w273;
 wire w274,w275,w276,w277,w278,w279,w280,w281;
 wire w282,w283,w284,w285,w286,w287,w288,w289;
 wire w290,w291,w292,w293,w294,w295,w296,w297;
 wire w298,w299,w300,w301,w302,w303,w304,w305;
 wire w306,w307,w308,w309,w310,w311,w312,w313;
 wire w314,w315,w316,w317,w318,w319,w320,w321;
 wire w322,w323,w324,w325,w326,w327,w328,w329;
 wire w330,w331,w332,w333,w334,w335,w336,w337;
 wire w338,w339,w340,w341,w342,w343,w344,w345;
 wire w346,w347,w348,w349,w350,w351,w352,w353;
 wire w354,w355,w356,w357,w358,w359,w360,w361;
 wire w362,w363,w364,w365,w366,w367,w368,w369;
 wire w370,w371,w372,w373,w374,w375,w376,w377;
 wire w378,w379,w380,w381,w382,w383,w384,w385;
 wire w386,w387,w388,w389,w390,w391,w392,w393;
 wire w394,w395,w396,w397,w398,w399,w400,w401;
 wire w402,w403,w404,w405,w406,w407,w408,w409;
 wire w410,w411,w412,w413,w414,w415,w416,w417;
 wire w418,w419,w420,w421,w422,w423,w424,w425;
 wire w426,w427,w428,w429,w430,w431,w432,w433;
 wire w434,w435,w436,w437,w438,w439,w440,w441;
 wire w442,w443,w444,w445,w446,w447,w448,w449;
 wire w450,w451,w452,w453,w454,w455,w456,w457;
 wire w458,w459,w460,w461,w462,w463,w464,w465;
 wire w466,w467,w468,w469,w470,w471,w472,w473;
 wire w474,w475,w476,w477,w478,w479,w480,w481;
 wire w482,w483,w484,w485,w486,w487,w488,w489;
 wire w490,w491,w492,w493,w494,w495,w496,w497;
 wire w498,w499,w500,w501,w502,w503,w504,w505;
 wire w506,w507,w508,w509,w510,w511,w512,w513;
 not #(2) NOT_1_1_1(w38,MC3);
 not #(8) NOT_2_2_2(w20,w38);
 pmos #(2) pmos_1_3_3_3(w38,vdd,MC3); //  
 nmos #(2) nmos_2_4_4_4(w38,vss,MC3); //  
 pmos #(8) pmos_1_5_5_5(w20,vdd,w38); //  
 nmos #(8) nmos_2_6_6_6(w20,vss,w38); //  
 pmos #(1) pmos_1_7_7(w40,vdd,w39); //  
 nmos #(2) nmos_2_8_8(w41,vss,w39); //  
 nmos #(2) nmos_3_9_9(w41,vss,w42); //  
 pmos #(2) pmos_4_10_10(w41,w40,w42); //  
 nmos #(3) nmos_5_11_11(w18,vss,w41); //  
 pmos #(3) pmos_6_12_12(w18,vdd,w41); //  
 pmos #(1) pmos_1_13_13(w43,vdd,MC2); //  
 nmos #(1) nmos_2_14_14(w43,vss,MC2); //  
 pmos #(1) pmos_1_1_15_15(w45,vdd,w44); //  
 nmos #(2) nmos_2_2_16_16(w46,vss,w44); //  
 nmos #(2) nmos_3_3_17_17(w46,vss,w47); //  
 pmos #(2) pmos_4_4_18_18(w46,w45,w47); //  
 nmos #(3) nmos_5_5_19_19(w19,vss,w46); //  
 pmos #(3) pmos_6_6_20_20(w19,vdd,w46); //  
 pmos #(1) pmos_1_7_21_21(w48,vdd,MC2); //  
 nmos #(1) nmos_2_8_22_22(w48,vss,MC2); //  
 nmos #(1) nmos_1_9_23_23(w49,vss,w48); //  
 pmos #(2) pmos_2_10_24_24(w50,vdd,MC1); //  
 pmos #(2) pmos_3_11_25_25(w50,vdd,w48); //  
 nmos #(2) nmos_4_12_26_26(w50,w49,MC1); //  
 nmos #(1) nmos_5_13_27_27(w44,vss,w50); //  
 pmos #(1) pmos_6_14_28_28(w44,vdd,w50); //  
 pmos #(1) pmos_1_15_29_29(w51,vdd,MC1); //  
 nmos #(1) nmos_2_16_30_30(w51,vss,MC1); //  
 nmos #(1) nmos_1_17_31_31(w52,vss,w51); //  
 pmos #(2) pmos_2_18_32_32(w53,vdd,MC2); //  
 pmos #(2) pmos_3_19_33_33(w53,vdd,w51); //  
 nmos #(2) nmos_4_20_34_34(w53,w52,MC2); //  
 nmos #(1) nmos_5_21_35_35(w47,vss,w53); //  
 pmos #(1) pmos_6_22_36_36(w47,vdd,w53); //  
 pmos #(1) pmos_1_37_37(w54,vdd,MC1); //  
 nmos #(1) nmos_2_38_38(w54,vss,MC1); //  
 nmos #(1) nmos_1_39_39(w55,vss,MC2); //  
 pmos #(2) pmos_2_40_40(w56,vdd,MC1); //  
 pmos #(2) pmos_3_41_41(w56,vdd,MC2); //  
 nmos #(2) nmos_4_42_42(w56,w55,MC1); //  
 nmos #(1) nmos_5_43_43(w57,vss,w56); //  
 pmos #(1) pmos_6_44_44(w57,vdd,w56); //  
 nmos #(1) nmos_1_45_45(w58,vss,MC3); //  
 pmos #(2) pmos_2_46_46(w60,vdd,w59); //  
 pmos #(2) pmos_3_47_47(w60,vdd,MC3); //  
 nmos #(2) nmos_4_48_48(w60,w58,w59); //  
 nmos #(1) nmos_5_49_49(w39,vss,w60); //  
 pmos #(1) pmos_6_50_50(w39,vdd,w60); //  
 nmos #(1) nmos_1_51_51(w61,vss,w43); //  
 pmos #(2) pmos_2_52_52(w62,vdd,w54); //  
 pmos #(2) pmos_3_53_53(w62,vdd,w43); //  
 nmos #(2) nmos_4_54_54(w62,w61,w54); //  
 nmos #(1) nmos_5_55_55(w59,vss,w62); //  
 pmos #(1) pmos_6_56_56(w59,vdd,w62); //  
 pmos #(1) pmos_1_57_57(w63,vdd,MC3); //  
 nmos #(1) nmos_2_58_58(w63,vss,MC3); //  
 nmos #(1) nmos_1_59_59(w64,vss,w63); //  
 pmos #(2) pmos_2_60_60(w65,vdd,w57); //  
 pmos #(2) pmos_3_61_61(w65,vdd,w63); //  
 nmos #(2) nmos_4_62_62(w65,w64,w57); //  
 nmos #(1) nmos_5_63_63(w42,vss,w65); //  
 pmos #(1) pmos_6_64_64(w42,vdd,w65); //  
 pmos #(1) pmos_1_1_1_65(w67,vdd,w66); //  
 nmos #(2) nmos_2_2_2_66(w68,vss,w66); //  
 nmos #(2) nmos_3_3_3_67(w68,vss,w69); //  
 pmos #(2) pmos_4_4_4_68(w68,w67,w69); //  
 nmos #(2) nmos_5_5_5_69(w70,vss,w68); //  
 pmos #(2) pmos_6_6_6_70(w70,vdd,w68); //  
 pmos #(1) pmos_1_1_7_7_71(w72,vdd,w71); //  
 nmos #(2) nmos_2_2_8_8_72(w73,vss,w71); //  
 nmos #(2) nmos_3_3_9_9_73(w73,vss,w74); //  
 pmos #(2) pmos_4_4_10_10_74(w73,w72,w74); //  
 nmos #(6) nmos_5_5_11_11_75(w24,vss,w73); //  
 pmos #(6) pmos_6_6_12_12_76(w24,vdd,w73); //  
 pmos #(1) pmos_1_7_13_13_77(w75,vdd,w23); //  
 nmos #(1) nmos_2_8_14_14_78(w75,vss,w23); //  
 nmos #(1) nmos_1_9_15_15_79(w76,vss,w75); //  
 pmos #(2) pmos_2_10_16_16_80(w77,vdd,w70); //  
 pmos #(2) pmos_3_11_17_17_81(w77,vdd,w75); //  
 nmos #(2) nmos_4_12_18_18_82(w77,w76,w70); //  
 nmos #(1) nmos_5_13_19_19_83(w71,vss,w77); //  
 pmos #(1) pmos_6_14_20_20_84(w71,vdd,w77); //  
 pmos #(1) pmos_1_15_21_21_85(w78,vdd,w70); //  
 nmos #(1) nmos_2_16_22_22_86(w78,vss,w70); //  
 nmos #(1) nmos_1_17_23_23_87(w79,vss,w78); //  
 pmos #(2) pmos_2_18_24_24_88(w80,vdd,w23); //  
 pmos #(2) pmos_3_19_25_25_89(w80,vdd,w78); //  
 nmos #(2) nmos_4_20_26_26_90(w80,w79,w23); //  
 nmos #(1) nmos_5_21_27_27_91(w74,vss,w80); //  
 pmos #(1) pmos_6_22_28_28_92(w74,vdd,w80); //  
 nmos #(1) nmos_1_29_29_93(w81,vss,w22); //  
 pmos #(2) pmos_2_30_30_94(w82,vdd,MP2); //  
 pmos #(2) pmos_3_31_31_95(w82,vdd,w22); //  
 nmos #(2) nmos_4_32_32_96(w82,w81,MP2); //  
 nmos #(1) nmos_5_33_33_97(w66,vss,w82); //  
 pmos #(1) pmos_6_34_34_98(w66,vdd,w82); //  
 nmos #(1) nmos_1_35_35_99(w83,vss,w21); //  
 pmos #(2) pmos_2_36_36_100(w84,vdd,MP3); //  
 pmos #(2) pmos_3_37_37_101(w84,vdd,w21); //  
 nmos #(2) nmos_4_38_38_102(w84,w83,MP3); //  
 nmos #(1) nmos_5_39_39_103(w69,vss,w84); //  
 pmos #(1) pmos_6_40_40_104(w69,vdd,w84); //  
 pmos #(1) pmos_1_1_41_105(w86,vdd,w85); //  
 nmos #(2) nmos_2_2_42_106(w87,vss,w85); //  
 nmos #(2) nmos_3_3_43_107(w87,vss,w88); //  
 pmos #(2) pmos_4_4_44_108(w87,w86,w88); //  
 nmos #(2) nmos_5_5_45_109(w89,vss,w87); //  
 pmos #(2) pmos_6_6_46_110(w89,vdd,w87); //  
 pmos #(1) pmos_1_1_7_47_111(w91,vdd,w90); //  
 nmos #(2) nmos_2_2_8_48_112(w92,vss,w90); //  
 nmos #(2) nmos_3_3_9_49_113(w92,vss,w93); //  
 pmos #(2) pmos_4_4_10_50_114(w92,w91,w93); //  
 nmos #(3) nmos_5_5_11_51_115(w27,vss,w92); //  
 pmos #(3) pmos_6_6_12_52_116(w27,vdd,w92); //  
 pmos #(1) pmos_1_7_13_53_117(w94,vdd,w23); //  
 nmos #(1) nmos_2_8_14_54_118(w94,vss,w23); //  
 nmos #(1) nmos_1_9_15_55_119(w95,vss,w94); //  
 pmos #(2) pmos_2_10_16_56_120(w96,vdd,w89); //  
 pmos #(2) pmos_3_11_17_57_121(w96,vdd,w94); //  
 nmos #(2) nmos_4_12_18_58_122(w96,w95,w89); //  
 nmos #(1) nmos_5_13_19_59_123(w90,vss,w96); //  
 pmos #(1) pmos_6_14_20_60_124(w90,vdd,w96); //  
 pmos #(1) pmos_1_15_21_61_125(w97,vdd,w89); //  
 nmos #(1) nmos_2_16_22_62_126(w97,vss,w89); //  
 nmos #(1) nmos_1_17_23_63_127(w98,vss,w97); //  
 pmos #(2) pmos_2_18_24_64_128(w99,vdd,w23); //  
 pmos #(2) pmos_3_19_25_65_129(w99,vdd,w97); //  
 nmos #(2) nmos_4_20_26_66_130(w99,w98,w23); //  
 nmos #(1) nmos_5_21_27_67_131(w93,vss,w99); //  
 pmos #(1) pmos_6_22_28_68_132(w93,vdd,w99); //  
 nmos #(1) nmos_1_29_69_133(w100,vss,w22); //  
 pmos #(2) pmos_2_30_70_134(w101,vdd,MP1); //  
 pmos #(2) pmos_3_31_71_135(w101,vdd,w22); //  
 nmos #(2) nmos_4_32_72_136(w101,w100,MP1); //  
 nmos #(1) nmos_5_33_73_137(w85,vss,w101); //  
 pmos #(1) pmos_6_34_74_138(w85,vdd,w101); //  
 nmos #(1) nmos_1_35_75_139(w102,vss,w21); //  
 pmos #(2) pmos_2_36_76_140(w103,vdd,MP2); //  
 pmos #(2) pmos_3_37_77_141(w103,vdd,w21); //  
 nmos #(2) nmos_4_38_78_142(w103,w102,MP2); //  
 nmos #(1) nmos_5_39_79_143(w88,vss,w103); //  
 pmos #(1) pmos_6_40_80_144(w88,vdd,w103); //  
 pmos #(1) pmos_1_1_81_145(w105,vdd,w104); //  
 nmos #(2) nmos_2_2_82_146(w106,vss,w104); //  
 nmos #(2) nmos_3_3_83_147(w106,vss,w107); //  
 pmos #(2) pmos_4_4_84_148(w106,w105,w107); //  
 nmos #(2) nmos_5_5_85_149(w108,vss,w106); //  
 pmos #(2) pmos_6_6_86_150(w108,vdd,w106); //  
 pmos #(1) pmos_1_1_7_87_151(w110,vdd,w109); //  
 nmos #(2) nmos_2_2_8_88_152(w111,vss,w109); //  
 nmos #(2) nmos_3_3_9_89_153(w111,vss,w112); //  
 pmos #(2) pmos_4_4_10_90_154(w111,w110,w112); //  
 nmos #(3) nmos_5_5_11_91_155(w25,vss,w111); //  
 pmos #(3) pmos_6_6_12_92_156(w25,vdd,w111); //  
 pmos #(1) pmos_1_7_13_93_157(w113,vdd,w23); //  
 nmos #(1) nmos_2_8_14_94_158(w113,vss,w23); //  
 nmos #(1) nmos_1_9_15_95_159(w114,vss,w113); //  
 pmos #(2) pmos_2_10_16_96_160(w115,vdd,w108); //  
 pmos #(2) pmos_3_11_17_97_161(w115,vdd,w113); //  
 nmos #(2) nmos_4_12_18_98_162(w115,w114,w108); //  
 nmos #(1) nmos_5_13_19_99_163(w109,vss,w115); //  
 pmos #(1) pmos_6_14_20_100_164(w109,vdd,w115); //  
 pmos #(1) pmos_1_15_21_101_165(w116,vdd,w108); //  
 nmos #(1) nmos_2_16_22_102_166(w116,vss,w108); //  
 nmos #(1) nmos_1_17_23_103_167(w117,vss,w116); //  
 pmos #(2) pmos_2_18_24_104_168(w118,vdd,w23); //  
 pmos #(2) pmos_3_19_25_105_169(w118,vdd,w116); //  
 nmos #(2) nmos_4_20_26_106_170(w118,w117,w23); //  
 nmos #(1) nmos_5_21_27_107_171(w112,vss,w118); //  
 pmos #(1) pmos_6_22_28_108_172(w112,vdd,w118); //  
 nmos #(1) nmos_1_29_109_173(w119,vss,w22); //  
 pmos #(2) pmos_2_30_110_174(w120,vdd,MP0); //  
 pmos #(2) pmos_3_31_111_175(w120,vdd,w22); //  
 nmos #(2) nmos_4_32_112_176(w120,w119,MP0); //  
 nmos #(1) nmos_5_33_113_177(w104,vss,w120); //  
 pmos #(1) pmos_6_34_114_178(w104,vdd,w120); //  
 nmos #(1) nmos_1_35_115_179(w121,vss,w21); //  
 pmos #(2) pmos_2_36_116_180(w122,vdd,MP1); //  
 pmos #(2) pmos_3_37_117_181(w122,vdd,w21); //  
 nmos #(2) nmos_4_38_118_182(w122,w121,MP1); //  
 nmos #(1) nmos_5_39_119_183(w107,vss,w122); //  
 pmos #(1) pmos_6_40_120_184(w107,vdd,w122); //  
 pmos #(1) pmos_1_1_121_185(w124,vdd,w123); //  
 nmos #(2) nmos_2_2_122_186(w125,vss,w123); //  
 nmos #(2) nmos_3_3_123_187(w125,vss,w126); //  
 pmos #(2) pmos_4_4_124_188(w125,w124,w126); //  
 nmos #(2) nmos_5_5_125_189(w127,vss,w125); //  
 pmos #(2) pmos_6_6_126_190(w127,vdd,w125); //  
 pmos #(1) pmos_1_1_7_127_191(w129,vdd,w128); //  
 nmos #(2) nmos_2_2_8_128_192(w130,vss,w128); //  
 nmos #(2) nmos_3_3_9_129_193(w130,vss,w131); //  
 pmos #(2) pmos_4_4_10_130_194(w130,w129,w131); //  
 nmos #(3) nmos_5_5_11_131_195(w26,vss,w130); //  
 pmos #(3) pmos_6_6_12_132_196(w26,vdd,w130); //  
 pmos #(1) pmos_1_7_13_133_197(w132,vdd,w23); //  
 nmos #(1) nmos_2_8_14_134_198(w132,vss,w23); //  
 nmos #(1) nmos_1_9_15_135_199(w133,vss,w132); //  
 pmos #(2) pmos_2_10_16_136_200(w134,vdd,w127); //  
 pmos #(2) pmos_3_11_17_137_201(w134,vdd,w132); //  
 nmos #(2) nmos_4_12_18_138_202(w134,w133,w127); //  
 nmos #(1) nmos_5_13_19_139_203(w128,vss,w134); //  
 pmos #(1) pmos_6_14_20_140_204(w128,vdd,w134); //  
 pmos #(1) pmos_1_15_21_141_205(w135,vdd,w127); //  
 nmos #(1) nmos_2_16_22_142_206(w135,vss,w127); //  
 nmos #(1) nmos_1_17_23_143_207(w136,vss,w135); //  
 pmos #(2) pmos_2_18_24_144_208(w137,vdd,w23); //  
 pmos #(2) pmos_3_19_25_145_209(w137,vdd,w135); //  
 nmos #(2) nmos_4_20_26_146_210(w137,w136,w23); //  
 nmos #(1) nmos_5_21_27_147_211(w131,vss,w137); //  
 pmos #(1) pmos_6_22_28_148_212(w131,vdd,w137); //  
 nmos #(1) nmos_1_29_149_213(w138,vss,w22); //  
 pmos #(2) pmos_2_30_150_214(w139,vdd,vss); //  
 pmos #(2) pmos_3_31_151_215(w139,vdd,w22); //  
 nmos #(2) nmos_4_32_152_216(w139,w138,vss); //  
 nmos #(1) nmos_5_33_153_217(w123,vss,w139); //  
 pmos #(1) pmos_6_34_154_218(w123,vdd,w139); //  
 nmos #(1) nmos_1_35_155_219(w140,vss,w21); //  
 pmos #(2) pmos_2_36_156_220(w141,vdd,MP0); //  
 pmos #(2) pmos_3_37_157_221(w141,vdd,w21); //  
 nmos #(2) nmos_4_38_158_222(w141,w140,MP0); //  
 nmos #(1) nmos_5_39_159_223(w126,vss,w141); //  
 pmos #(1) pmos_6_40_160_224(w126,vdd,w141); //  
 pmos #(1) pmos_1_1_1_225(w143,vdd,w142); //  
 nmos #(2) nmos_2_2_2_226(w144,vss,w142); //  
 nmos #(2) nmos_3_3_3_227(w144,vss,w145); //  
 pmos #(2) pmos_4_4_4_228(w144,w143,w145); //  
 nmos #(2) nmos_5_5_5_229(w146,vss,w144); //  
 pmos #(2) pmos_6_6_6_230(w146,vdd,w144); //  
 pmos #(1) pmos_1_1_7_7_231(w148,vdd,w147); //  
 nmos #(2) nmos_2_2_8_8_232(w149,vss,w147); //  
 nmos #(2) nmos_3_3_9_9_233(w149,vss,w150); //  
 pmos #(2) pmos_4_4_10_10_234(w149,w148,w150); //  
 nmos #(6) nmos_5_5_11_11_235(w28,vss,w149); //  
 pmos #(6) pmos_6_6_12_12_236(w28,vdd,w149); //  
 pmos #(1) pmos_1_7_13_13_237(w151,vdd,w20); //  
 nmos #(1) nmos_2_8_14_14_238(w151,vss,w20); //  
 nmos #(1) nmos_1_9_15_15_239(w152,vss,w151); //  
 pmos #(2) pmos_2_10_16_16_240(w153,vdd,w146); //  
 pmos #(2) pmos_3_11_17_17_241(w153,vdd,w151); //  
 nmos #(2) nmos_4_12_18_18_242(w153,w152,w146); //  
 nmos #(1) nmos_5_13_19_19_243(w147,vss,w153); //  
 pmos #(1) pmos_6_14_20_20_244(w147,vdd,w153); //  
 pmos #(1) pmos_1_15_21_21_245(w154,vdd,w146); //  
 nmos #(1) nmos_2_16_22_22_246(w154,vss,w146); //  
 nmos #(1) nmos_1_17_23_23_247(w155,vss,w154); //  
 pmos #(2) pmos_2_18_24_24_248(w156,vdd,w20); //  
 pmos #(2) pmos_3_19_25_25_249(w156,vdd,w154); //  
 nmos #(2) nmos_4_20_26_26_250(w156,w155,w20); //  
 nmos #(1) nmos_5_21_27_27_251(w150,vss,w156); //  
 pmos #(1) pmos_6_22_28_28_252(w150,vdd,w156); //  
 nmos #(1) nmos_1_29_29_253(w157,vss,w18); //  
 pmos #(2) pmos_2_30_30_254(w158,vdd,MP2); //  
 pmos #(2) pmos_3_31_31_255(w158,vdd,w18); //  
 nmos #(2) nmos_4_32_32_256(w158,w157,MP2); //  
 nmos #(1) nmos_5_33_33_257(w142,vss,w158); //  
 pmos #(1) pmos_6_34_34_258(w142,vdd,w158); //  
 nmos #(1) nmos_1_35_35_259(w159,vss,w19); //  
 pmos #(2) pmos_2_36_36_260(w160,vdd,MP3); //  
 pmos #(2) pmos_3_37_37_261(w160,vdd,w19); //  
 nmos #(2) nmos_4_38_38_262(w160,w159,MP3); //  
 nmos #(1) nmos_5_39_39_263(w145,vss,w160); //  
 pmos #(1) pmos_6_40_40_264(w145,vdd,w160); //  
 pmos #(1) pmos_1_1_41_265(w162,vdd,w161); //  
 nmos #(2) nmos_2_2_42_266(w163,vss,w161); //  
 nmos #(2) nmos_3_3_43_267(w163,vss,w164); //  
 pmos #(2) pmos_4_4_44_268(w163,w162,w164); //  
 nmos #(2) nmos_5_5_45_269(w165,vss,w163); //  
 pmos #(2) pmos_6_6_46_270(w165,vdd,w163); //  
 pmos #(1) pmos_1_1_7_47_271(w167,vdd,w166); //  
 nmos #(2) nmos_2_2_8_48_272(w168,vss,w166); //  
 nmos #(2) nmos_3_3_9_49_273(w168,vss,w169); //  
 pmos #(2) pmos_4_4_10_50_274(w168,w167,w169); //  
 nmos #(3) nmos_5_5_11_51_275(w31,vss,w168); //  
 pmos #(3) pmos_6_6_12_52_276(w31,vdd,w168); //  
 pmos #(1) pmos_1_7_13_53_277(w170,vdd,w20); //  
 nmos #(1) nmos_2_8_14_54_278(w170,vss,w20); //  
 nmos #(1) nmos_1_9_15_55_279(w171,vss,w170); //  
 pmos #(2) pmos_2_10_16_56_280(w172,vdd,w165); //  
 pmos #(2) pmos_3_11_17_57_281(w172,vdd,w170); //  
 nmos #(2) nmos_4_12_18_58_282(w172,w171,w165); //  
 nmos #(1) nmos_5_13_19_59_283(w166,vss,w172); //  
 pmos #(1) pmos_6_14_20_60_284(w166,vdd,w172); //  
 pmos #(1) pmos_1_15_21_61_285(w173,vdd,w165); //  
 nmos #(1) nmos_2_16_22_62_286(w173,vss,w165); //  
 nmos #(1) nmos_1_17_23_63_287(w174,vss,w173); //  
 pmos #(2) pmos_2_18_24_64_288(w175,vdd,w20); //  
 pmos #(2) pmos_3_19_25_65_289(w175,vdd,w173); //  
 nmos #(2) nmos_4_20_26_66_290(w175,w174,w20); //  
 nmos #(1) nmos_5_21_27_67_291(w169,vss,w175); //  
 pmos #(1) pmos_6_22_28_68_292(w169,vdd,w175); //  
 nmos #(1) nmos_1_29_69_293(w176,vss,w18); //  
 pmos #(2) pmos_2_30_70_294(w177,vdd,MP1); //  
 pmos #(2) pmos_3_31_71_295(w177,vdd,w18); //  
 nmos #(2) nmos_4_32_72_296(w177,w176,MP1); //  
 nmos #(1) nmos_5_33_73_297(w161,vss,w177); //  
 pmos #(1) pmos_6_34_74_298(w161,vdd,w177); //  
 nmos #(1) nmos_1_35_75_299(w178,vss,w19); //  
 pmos #(2) pmos_2_36_76_300(w179,vdd,MP2); //  
 pmos #(2) pmos_3_37_77_301(w179,vdd,w19); //  
 nmos #(2) nmos_4_38_78_302(w179,w178,MP2); //  
 nmos #(1) nmos_5_39_79_303(w164,vss,w179); //  
 pmos #(1) pmos_6_40_80_304(w164,vdd,w179); //  
 pmos #(1) pmos_1_1_81_305(w181,vdd,w180); //  
 nmos #(2) nmos_2_2_82_306(w182,vss,w180); //  
 nmos #(2) nmos_3_3_83_307(w182,vss,w183); //  
 pmos #(2) pmos_4_4_84_308(w182,w181,w183); //  
 nmos #(2) nmos_5_5_85_309(w184,vss,w182); //  
 pmos #(2) pmos_6_6_86_310(w184,vdd,w182); //  
 pmos #(1) pmos_1_1_7_87_311(w186,vdd,w185); //  
 nmos #(2) nmos_2_2_8_88_312(w187,vss,w185); //  
 nmos #(2) nmos_3_3_9_89_313(w187,vss,w188); //  
 pmos #(2) pmos_4_4_10_90_314(w187,w186,w188); //  
 nmos #(3) nmos_5_5_11_91_315(w29,vss,w187); //  
 pmos #(3) pmos_6_6_12_92_316(w29,vdd,w187); //  
 pmos #(1) pmos_1_7_13_93_317(w189,vdd,w20); //  
 nmos #(1) nmos_2_8_14_94_318(w189,vss,w20); //  
 nmos #(1) nmos_1_9_15_95_319(w190,vss,w189); //  
 pmos #(2) pmos_2_10_16_96_320(w191,vdd,w184); //  
 pmos #(2) pmos_3_11_17_97_321(w191,vdd,w189); //  
 nmos #(2) nmos_4_12_18_98_322(w191,w190,w184); //  
 nmos #(1) nmos_5_13_19_99_323(w185,vss,w191); //  
 pmos #(1) pmos_6_14_20_100_324(w185,vdd,w191); //  
 pmos #(1) pmos_1_15_21_101_325(w192,vdd,w184); //  
 nmos #(1) nmos_2_16_22_102_326(w192,vss,w184); //  
 nmos #(1) nmos_1_17_23_103_327(w193,vss,w192); //  
 pmos #(2) pmos_2_18_24_104_328(w194,vdd,w20); //  
 pmos #(2) pmos_3_19_25_105_329(w194,vdd,w192); //  
 nmos #(2) nmos_4_20_26_106_330(w194,w193,w20); //  
 nmos #(1) nmos_5_21_27_107_331(w188,vss,w194); //  
 pmos #(1) pmos_6_22_28_108_332(w188,vdd,w194); //  
 nmos #(1) nmos_1_29_109_333(w195,vss,w18); //  
 pmos #(2) pmos_2_30_110_334(w196,vdd,MP0); //  
 pmos #(2) pmos_3_31_111_335(w196,vdd,w18); //  
 nmos #(2) nmos_4_32_112_336(w196,w195,MP0); //  
 nmos #(1) nmos_5_33_113_337(w180,vss,w196); //  
 pmos #(1) pmos_6_34_114_338(w180,vdd,w196); //  
 nmos #(1) nmos_1_35_115_339(w197,vss,w19); //  
 pmos #(2) pmos_2_36_116_340(w198,vdd,MP1); //  
 pmos #(2) pmos_3_37_117_341(w198,vdd,w19); //  
 nmos #(2) nmos_4_38_118_342(w198,w197,MP1); //  
 nmos #(1) nmos_5_39_119_343(w183,vss,w198); //  
 pmos #(1) pmos_6_40_120_344(w183,vdd,w198); //  
 pmos #(1) pmos_1_1_121_345(w200,vdd,w199); //  
 nmos #(2) nmos_2_2_122_346(w201,vss,w199); //  
 nmos #(2) nmos_3_3_123_347(w201,vss,w202); //  
 pmos #(2) pmos_4_4_124_348(w201,w200,w202); //  
 nmos #(2) nmos_5_5_125_349(w203,vss,w201); //  
 pmos #(2) pmos_6_6_126_350(w203,vdd,w201); //  
 pmos #(1) pmos_1_1_7_127_351(w205,vdd,w204); //  
 nmos #(2) nmos_2_2_8_128_352(w206,vss,w204); //  
 nmos #(2) nmos_3_3_9_129_353(w206,vss,w207); //  
 pmos #(2) pmos_4_4_10_130_354(w206,w205,w207); //  
 nmos #(3) nmos_5_5_11_131_355(w30,vss,w206); //  
 pmos #(3) pmos_6_6_12_132_356(w30,vdd,w206); //  
 pmos #(1) pmos_1_7_13_133_357(w208,vdd,w20); //  
 nmos #(1) nmos_2_8_14_134_358(w208,vss,w20); //  
 nmos #(1) nmos_1_9_15_135_359(w209,vss,w208); //  
 pmos #(2) pmos_2_10_16_136_360(w210,vdd,w203); //  
 pmos #(2) pmos_3_11_17_137_361(w210,vdd,w208); //  
 nmos #(2) nmos_4_12_18_138_362(w210,w209,w203); //  
 nmos #(1) nmos_5_13_19_139_363(w204,vss,w210); //  
 pmos #(1) pmos_6_14_20_140_364(w204,vdd,w210); //  
 pmos #(1) pmos_1_15_21_141_365(w211,vdd,w203); //  
 nmos #(1) nmos_2_16_22_142_366(w211,vss,w203); //  
 nmos #(1) nmos_1_17_23_143_367(w212,vss,w211); //  
 pmos #(2) pmos_2_18_24_144_368(w213,vdd,w20); //  
 pmos #(2) pmos_3_19_25_145_369(w213,vdd,w211); //  
 nmos #(2) nmos_4_20_26_146_370(w213,w212,w20); //  
 nmos #(1) nmos_5_21_27_147_371(w207,vss,w213); //  
 pmos #(1) pmos_6_22_28_148_372(w207,vdd,w213); //  
 nmos #(1) nmos_1_29_149_373(w214,vss,w18); //  
 pmos #(2) pmos_2_30_150_374(w215,vdd,vss); //  
 pmos #(2) pmos_3_31_151_375(w215,vdd,w18); //  
 nmos #(2) nmos_4_32_152_376(w215,w214,vss); //  
 nmos #(1) nmos_5_33_153_377(w199,vss,w215); //  
 pmos #(1) pmos_6_34_154_378(w199,vdd,w215); //  
 nmos #(1) nmos_1_35_155_379(w216,vss,w19); //  
 pmos #(2) pmos_2_36_156_380(w217,vdd,MP0); //  
 pmos #(2) pmos_3_37_157_381(w217,vdd,w19); //  
 nmos #(2) nmos_4_38_158_382(w217,w216,MP0); //  
 nmos #(1) nmos_5_39_159_383(w202,vss,w217); //  
 pmos #(1) pmos_6_40_160_384(w202,vdd,w217); //  
 pmos #(1) pmos_1_1_1_1_1_385(w219,vdd,w218); //  
 nmos #(2) nmos_2_2_2_2_2_386(w220,vss,w218); //  
 nmos #(2) nmos_3_3_3_3_3_387(w220,vss,w221); //  
 pmos #(2) pmos_4_4_4_4_4_388(w220,w219,w221); //  
 nmos #(3) nmos_5_5_5_5_5_389(w35,vss,w220); //  
 pmos #(3) pmos_6_6_6_6_6_390(w35,vdd,w220); //  
 pmos #(1) pmos_1_7_7_7_7_391(w223,vdd,w222); //  
 nmos #(1) nmos_2_8_8_8_8_392(w223,vss,w222); //  
 nmos #(1) nmos_1_9_9_9_9_393(w224,vss,w223); //  
 pmos #(2) pmos_2_10_10_10_10_394(w226,vdd,w225); //  
 pmos #(2) pmos_3_11_11_11_11_395(w226,vdd,w223); //  
 nmos #(2) nmos_4_12_12_12_12_396(w226,w224,w225); //  
 nmos #(1) nmos_5_13_13_13_13_397(w218,vss,w226); //  
 pmos #(1) pmos_6_14_14_14_14_398(w218,vdd,w226); //  
 pmos #(1) pmos_1_15_15_15_15_399(w227,vdd,w225); //  
 nmos #(1) nmos_2_16_16_16_16_400(w227,vss,w225); //  
 nmos #(1) nmos_1_17_17_17_17_401(w228,vss,w227); //  
 pmos #(2) pmos_2_18_18_18_18_402(w229,vdd,w222); //  
 pmos #(2) pmos_3_19_19_19_19_403(w229,vdd,w227); //  
 nmos #(2) nmos_4_20_20_20_20_404(w229,w228,w222); //  
 nmos #(1) nmos_5_21_21_21_21_405(w221,vss,w229); //  
 pmos #(1) pmos_6_22_22_22_22_406(w221,vdd,w229); //  
 nmos #(1) nmos_1_23_23_23_407(w230,vss,w225); //  
 pmos #(2) pmos_2_24_24_24_408(w231,vdd,w222); //  
 pmos #(2) pmos_3_25_25_25_409(w231,vdd,w225); //  
 nmos #(2) nmos_4_26_26_26_410(w231,w230,w222); //  
 nmos #(1) nmos_5_27_27_27_411(w232,vss,w231); //  
 pmos #(1) pmos_6_28_28_28_412(w232,vdd,w231); //  
 pmos #(1) pmos_1_1_1_29_29_413(w234,vdd,w233); //  
 nmos #(2) nmos_2_2_2_30_30_414(w235,vss,w233); //  
 nmos #(2) nmos_3_3_3_31_31_415(w235,vss,w236); //  
 pmos #(2) pmos_4_4_4_32_32_416(w235,w234,w236); //  
 nmos #(4) nmos_5_5_5_33_33_417(w222,vss,w235); //  
 pmos #(4) pmos_6_6_6_34_34_418(w222,vdd,w235); //  
 pmos #(1) pmos_1_7_7_35_35_419(w237,vdd,w24); //  
 nmos #(1) nmos_2_8_8_36_36_420(w237,vss,w24); //  
 nmos #(1) nmos_1_9_9_37_37_421(w238,vss,w237); //  
 pmos #(2) pmos_2_10_10_38_38_422(w239,vdd,vss); //  
 pmos #(2) pmos_3_11_11_39_39_423(w239,vdd,w237); //  
 nmos #(2) nmos_4_12_12_40_40_424(w239,w238,vss); //  
 nmos #(1) nmos_5_13_13_41_41_425(w233,vss,w239); //  
 pmos #(1) pmos_6_14_14_42_42_426(w233,vdd,w239); //  
 pmos #(1) pmos_1_15_15_43_43_427(w240,vdd,vss); //  
 nmos #(1) nmos_2_16_16_44_44_428(w240,vss,vss); //  
 nmos #(1) nmos_1_17_17_45_45_429(w241,vss,w240); //  
 pmos #(2) pmos_2_18_18_46_46_430(w242,vdd,w24); //  
 pmos #(2) pmos_3_19_19_47_47_431(w242,vdd,w240); //  
 nmos #(2) nmos_4_20_20_48_48_432(w242,w241,w24); //  
 nmos #(1) nmos_5_21_21_49_49_433(w236,vss,w242); //  
 pmos #(1) pmos_6_22_22_50_50_434(w236,vdd,w242); //  
 nmos #(1) nmos_1_23_51_51_435(w243,vss,vss); //  
 pmos #(2) pmos_2_24_52_52_436(w244,vdd,w24); //  
 pmos #(2) pmos_3_25_53_53_437(w244,vdd,vss); //  
 nmos #(2) nmos_4_26_54_54_438(w244,w243,w24); //  
 nmos #(1) nmos_5_27_55_55_439(w245,vss,w244); //  
 pmos #(1) pmos_6_28_56_56_440(w245,vdd,w244); //  
 pmos #(1) pmos_1_57_57_441(w246,vdd,w245); //  
 nmos #(2) nmos_2_58_58_442(w247,vss,w245); //  
 nmos #(2) nmos_3_59_59_443(w247,vss,w232); //  
 pmos #(2) pmos_4_60_60_444(w247,w246,w232); //  
 nmos #(4) nmos_5_61_61_445(w248,vss,w247); //  
 pmos #(4) pmos_6_62_62_446(w248,vdd,w247); //  
 pmos #(1) pmos_1_1_1_1_63_447(w250,vdd,w249); //  
 nmos #(2) nmos_2_2_2_2_64_448(w251,vss,w249); //  
 nmos #(2) nmos_3_3_3_3_65_449(w251,vss,w252); //  
 pmos #(2) pmos_4_4_4_4_66_450(w251,w250,w252); //  
 nmos #(1) nmos_5_5_5_5_67_451(PROD0,vss,w251); //  
 pmos #(1) pmos_6_6_6_6_68_452(PROD0,vdd,w251); //  
 pmos #(1) pmos_1_7_7_7_69_453(w254,vdd,w253); //  
 nmos #(1) nmos_2_8_8_8_70_454(w254,vss,w253); //  
 nmos #(1) nmos_1_9_9_9_71_455(w255,vss,w254); //  
 pmos #(2) pmos_2_10_10_10_72_456(w256,vdd,w23); //  
 pmos #(2) pmos_3_11_11_11_73_457(w256,vdd,w254); //  
 nmos #(2) nmos_4_12_12_12_74_458(w256,w255,w23); //  
 nmos #(1) nmos_5_13_13_13_75_459(w249,vss,w256); //  
 pmos #(1) pmos_6_14_14_14_76_460(w249,vdd,w256); //  
 pmos #(1) pmos_1_15_15_15_77_461(w257,vdd,w23); //  
 nmos #(1) nmos_2_16_16_16_78_462(w257,vss,w23); //  
 nmos #(1) nmos_1_17_17_17_79_463(w258,vss,w257); //  
 pmos #(2) pmos_2_18_18_18_80_464(w259,vdd,w253); //  
 pmos #(2) pmos_3_19_19_19_81_465(w259,vdd,w257); //  
 nmos #(2) nmos_4_20_20_20_82_466(w259,w258,w253); //  
 nmos #(1) nmos_5_21_21_21_83_467(w252,vss,w259); //  
 pmos #(1) pmos_6_22_22_22_84_468(w252,vdd,w259); //  
 nmos #(1) nmos_1_23_23_85_469(w260,vss,w23); //  
 pmos #(2) pmos_2_24_24_86_470(w261,vdd,w253); //  
 pmos #(2) pmos_3_25_25_87_471(w261,vdd,w23); //  
 nmos #(2) nmos_4_26_26_88_472(w261,w260,w253); //  
 nmos #(1) nmos_5_27_27_89_473(w262,vss,w261); //  
 pmos #(1) pmos_6_28_28_90_474(w262,vdd,w261); //  
 pmos #(1) pmos_1_1_1_29_91_475(w264,vdd,w263); //  
 nmos #(2) nmos_2_2_2_30_92_476(w265,vss,w263); //  
 nmos #(2) nmos_3_3_3_31_93_477(w265,vss,w266); //  
 pmos #(2) pmos_4_4_4_32_94_478(w265,w264,w266); //  
 nmos #(4) nmos_5_5_5_33_95_479(w253,vss,w265); //  
 pmos #(4) pmos_6_6_6_34_96_480(w253,vdd,w265); //  
 pmos #(1) pmos_1_7_7_35_97_481(w267,vdd,w26); //  
 nmos #(1) nmos_2_8_8_36_98_482(w267,vss,w26); //  
 nmos #(1) nmos_1_9_9_37_99_483(w268,vss,w267); //  
 pmos #(2) pmos_2_10_10_38_100_484(w269,vdd,vss); //  
 pmos #(2) pmos_3_11_11_39_101_485(w269,vdd,w267); //  
 nmos #(2) nmos_4_12_12_40_102_486(w269,w268,vss); //  
 nmos #(1) nmos_5_13_13_41_103_487(w263,vss,w269); //  
 pmos #(1) pmos_6_14_14_42_104_488(w263,vdd,w269); //  
 pmos #(1) pmos_1_15_15_43_105_489(w270,vdd,vss); //  
 nmos #(1) nmos_2_16_16_44_106_490(w270,vss,vss); //  
 nmos #(1) nmos_1_17_17_45_107_491(w271,vss,w270); //  
 pmos #(2) pmos_2_18_18_46_108_492(w272,vdd,w26); //  
 pmos #(2) pmos_3_19_19_47_109_493(w272,vdd,w270); //  
 nmos #(2) nmos_4_20_20_48_110_494(w272,w271,w26); //  
 nmos #(1) nmos_5_21_21_49_111_495(w266,vss,w272); //  
 pmos #(1) pmos_6_22_22_50_112_496(w266,vdd,w272); //  
 nmos #(1) nmos_1_23_51_113_497(w273,vss,vss); //  
 pmos #(2) pmos_2_24_52_114_498(w274,vdd,w26); //  
 pmos #(2) pmos_3_25_53_115_499(w274,vdd,vss); //  
 nmos #(2) nmos_4_26_54_116_500(w274,w273,w26); //  
 nmos #(1) nmos_5_27_55_117_501(w275,vss,w274); //  
 pmos #(1) pmos_6_28_56_118_502(w275,vdd,w274); //  
 pmos #(1) pmos_1_57_119_503(w276,vdd,w275); //  
 nmos #(2) nmos_2_58_120_504(w277,vss,w275); //  
 nmos #(2) nmos_3_59_121_505(w277,vss,w262); //  
 pmos #(2) pmos_4_60_122_506(w277,w276,w262); //  
 nmos #(4) nmos_5_61_123_507(w278,vss,w277); //  
 pmos #(4) pmos_6_62_124_508(w278,vdd,w277); //  
 pmos #(1) pmos_1_1_1_1_125_509(w280,vdd,w279); //  
 nmos #(2) nmos_2_2_2_2_126_510(w281,vss,w279); //  
 nmos #(2) nmos_3_3_3_3_127_511(w281,vss,w282); //  
 pmos #(2) pmos_4_4_4_4_128_512(w281,w280,w282); //  
 nmos #(1) nmos_5_5_5_5_129_513(PROD1,vss,w281); //  
 pmos #(1) pmos_6_6_6_6_130_514(PROD1,vdd,w281); //  
 pmos #(1) pmos_1_7_7_7_131_515(w284,vdd,w283); //  
 nmos #(1) nmos_2_8_8_8_132_516(w284,vss,w283); //  
 nmos #(1) nmos_1_9_9_9_133_517(w285,vss,w284); //  
 pmos #(2) pmos_2_10_10_10_134_518(w286,vdd,w278); //  
 pmos #(2) pmos_3_11_11_11_135_519(w286,vdd,w284); //  
 nmos #(2) nmos_4_12_12_12_136_520(w286,w285,w278); //  
 nmos #(1) nmos_5_13_13_13_137_521(w279,vss,w286); //  
 pmos #(1) pmos_6_14_14_14_138_522(w279,vdd,w286); //  
 pmos #(1) pmos_1_15_15_15_139_523(w287,vdd,w278); //  
 nmos #(1) nmos_2_16_16_16_140_524(w287,vss,w278); //  
 nmos #(1) nmos_1_17_17_17_141_525(w288,vss,w287); //  
 pmos #(2) pmos_2_18_18_18_142_526(w289,vdd,w283); //  
 pmos #(2) pmos_3_19_19_19_143_527(w289,vdd,w287); //  
 nmos #(2) nmos_4_20_20_20_144_528(w289,w288,w283); //  
 nmos #(1) nmos_5_21_21_21_145_529(w282,vss,w289); //  
 pmos #(1) pmos_6_22_22_22_146_530(w282,vdd,w289); //  
 nmos #(1) nmos_1_23_23_147_531(w290,vss,w278); //  
 pmos #(2) pmos_2_24_24_148_532(w291,vdd,w283); //  
 pmos #(2) pmos_3_25_25_149_533(w291,vdd,w278); //  
 nmos #(2) nmos_4_26_26_150_534(w291,w290,w283); //  
 nmos #(1) nmos_5_27_27_151_535(w292,vss,w291); //  
 pmos #(1) pmos_6_28_28_152_536(w292,vdd,w291); //  
 pmos #(1) pmos_1_1_1_29_153_537(w294,vdd,w293); //  
 nmos #(2) nmos_2_2_2_30_154_538(w295,vss,w293); //  
 nmos #(2) nmos_3_3_3_31_155_539(w295,vss,w296); //  
 pmos #(2) pmos_4_4_4_32_156_540(w295,w294,w296); //  
 nmos #(4) nmos_5_5_5_33_157_541(w283,vss,w295); //  
 pmos #(4) pmos_6_6_6_34_158_542(w283,vdd,w295); //  
 pmos #(1) pmos_1_7_7_35_159_543(w297,vdd,w25); //  
 nmos #(1) nmos_2_8_8_36_160_544(w297,vss,w25); //  
 nmos #(1) nmos_1_9_9_37_161_545(w298,vss,w297); //  
 pmos #(2) pmos_2_10_10_38_162_546(w299,vdd,vss); //  
 pmos #(2) pmos_3_11_11_39_163_547(w299,vdd,w297); //  
 nmos #(2) nmos_4_12_12_40_164_548(w299,w298,vss); //  
 nmos #(1) nmos_5_13_13_41_165_549(w293,vss,w299); //  
 pmos #(1) pmos_6_14_14_42_166_550(w293,vdd,w299); //  
 pmos #(1) pmos_1_15_15_43_167_551(w300,vdd,vss); //  
 nmos #(1) nmos_2_16_16_44_168_552(w300,vss,vss); //  
 nmos #(1) nmos_1_17_17_45_169_553(w301,vss,w300); //  
 pmos #(2) pmos_2_18_18_46_170_554(w302,vdd,w25); //  
 pmos #(2) pmos_3_19_19_47_171_555(w302,vdd,w300); //  
 nmos #(2) nmos_4_20_20_48_172_556(w302,w301,w25); //  
 nmos #(1) nmos_5_21_21_49_173_557(w296,vss,w302); //  
 pmos #(1) pmos_6_22_22_50_174_558(w296,vdd,w302); //  
 nmos #(1) nmos_1_23_51_175_559(w303,vss,vss); //  
 pmos #(2) pmos_2_24_52_176_560(w304,vdd,w25); //  
 pmos #(2) pmos_3_25_53_177_561(w304,vdd,vss); //  
 nmos #(2) nmos_4_26_54_178_562(w304,w303,w25); //  
 nmos #(1) nmos_5_27_55_179_563(w305,vss,w304); //  
 pmos #(1) pmos_6_28_56_180_564(w305,vdd,w304); //  
 pmos #(1) pmos_1_57_181_565(w306,vdd,w305); //  
 nmos #(2) nmos_2_58_182_566(w307,vss,w305); //  
 nmos #(2) nmos_3_59_183_567(w307,vss,w292); //  
 pmos #(2) pmos_4_60_184_568(w307,w306,w292); //  
 nmos #(4) nmos_5_61_185_569(w308,vss,w307); //  
 pmos #(4) pmos_6_62_186_570(w308,vdd,w307); //  
 pmos #(1) pmos_1_1_1_1_187_571(w310,vdd,w309); //  
 nmos #(2) nmos_2_2_2_2_188_572(w311,vss,w309); //  
 nmos #(2) nmos_3_3_3_3_189_573(w311,vss,w312); //  
 pmos #(2) pmos_4_4_4_4_190_574(w311,w310,w312); //  
 nmos #(3) nmos_5_5_5_5_191_575(w36,vss,w311); //  
 pmos #(3) pmos_6_6_6_6_192_576(w36,vdd,w311); //  
 pmos #(1) pmos_1_7_7_7_193_577(w314,vdd,w313); //  
 nmos #(1) nmos_2_8_8_8_194_578(w314,vss,w313); //  
 nmos #(1) nmos_1_9_9_9_195_579(w315,vss,w314); //  
 pmos #(2) pmos_2_10_10_10_196_580(w316,vdd,w308); //  
 pmos #(2) pmos_3_11_11_11_197_581(w316,vdd,w314); //  
 nmos #(2) nmos_4_12_12_12_198_582(w316,w315,w308); //  
 nmos #(1) nmos_5_13_13_13_199_583(w309,vss,w316); //  
 pmos #(1) pmos_6_14_14_14_200_584(w309,vdd,w316); //  
 pmos #(1) pmos_1_15_15_15_201_585(w317,vdd,w308); //  
 nmos #(1) nmos_2_16_16_16_202_586(w317,vss,w308); //  
 nmos #(1) nmos_1_17_17_17_203_587(w318,vss,w317); //  
 pmos #(2) pmos_2_18_18_18_204_588(w319,vdd,w313); //  
 pmos #(2) pmos_3_19_19_19_205_589(w319,vdd,w317); //  
 nmos #(2) nmos_4_20_20_20_206_590(w319,w318,w313); //  
 nmos #(1) nmos_5_21_21_21_207_591(w312,vss,w319); //  
 pmos #(1) pmos_6_22_22_22_208_592(w312,vdd,w319); //  
 nmos #(1) nmos_1_23_23_209_593(w320,vss,w308); //  
 pmos #(2) pmos_2_24_24_210_594(w321,vdd,w313); //  
 pmos #(2) pmos_3_25_25_211_595(w321,vdd,w308); //  
 nmos #(2) nmos_4_26_26_212_596(w321,w320,w313); //  
 nmos #(1) nmos_5_27_27_213_597(w322,vss,w321); //  
 pmos #(1) pmos_6_28_28_214_598(w322,vdd,w321); //  
 pmos #(1) pmos_1_1_1_29_215_599(w324,vdd,w323); //  
 nmos #(2) nmos_2_2_2_30_216_600(w325,vss,w323); //  
 nmos #(2) nmos_3_3_3_31_217_601(w325,vss,w326); //  
 pmos #(2) pmos_4_4_4_32_218_602(w325,w324,w326); //  
 nmos #(4) nmos_5_5_5_33_219_603(w313,vss,w325); //  
 pmos #(4) pmos_6_6_6_34_220_604(w313,vdd,w325); //  
 pmos #(1) pmos_1_7_7_35_221_605(w327,vdd,w27); //  
 nmos #(1) nmos_2_8_8_36_222_606(w327,vss,w27); //  
 nmos #(1) nmos_1_9_9_37_223_607(w328,vss,w327); //  
 pmos #(2) pmos_2_10_10_38_224_608(w329,vdd,vss); //  
 pmos #(2) pmos_3_11_11_39_225_609(w329,vdd,w327); //  
 nmos #(2) nmos_4_12_12_40_226_610(w329,w328,vss); //  
 nmos #(1) nmos_5_13_13_41_227_611(w323,vss,w329); //  
 pmos #(1) pmos_6_14_14_42_228_612(w323,vdd,w329); //  
 pmos #(1) pmos_1_15_15_43_229_613(w330,vdd,vss); //  
 nmos #(1) nmos_2_16_16_44_230_614(w330,vss,vss); //  
 nmos #(1) nmos_1_17_17_45_231_615(w331,vss,w330); //  
 pmos #(2) pmos_2_18_18_46_232_616(w332,vdd,w27); //  
 pmos #(2) pmos_3_19_19_47_233_617(w332,vdd,w330); //  
 nmos #(2) nmos_4_20_20_48_234_618(w332,w331,w27); //  
 nmos #(1) nmos_5_21_21_49_235_619(w326,vss,w332); //  
 pmos #(1) pmos_6_22_22_50_236_620(w326,vdd,w332); //  
 nmos #(1) nmos_1_23_51_237_621(w333,vss,vss); //  
 pmos #(2) pmos_2_24_52_238_622(w334,vdd,w27); //  
 pmos #(2) pmos_3_25_53_239_623(w334,vdd,vss); //  
 nmos #(2) nmos_4_26_54_240_624(w334,w333,w27); //  
 nmos #(1) nmos_5_27_55_241_625(w335,vss,w334); //  
 pmos #(1) pmos_6_28_56_242_626(w335,vdd,w334); //  
 pmos #(1) pmos_1_57_243_627(w336,vdd,w335); //  
 nmos #(2) nmos_2_58_244_628(w337,vss,w335); //  
 nmos #(2) nmos_3_59_245_629(w337,vss,w322); //  
 pmos #(2) pmos_4_60_246_630(w337,w336,w322); //  
 nmos #(4) nmos_5_61_247_631(w225,vss,w337); //  
 pmos #(4) pmos_6_62_248_632(w225,vdd,w337); //  
 pmos #(1) pmos_1_1_1_1_249_633(w339,vdd,w338); //  
 nmos #(2) nmos_2_2_2_2_250_634(w340,vss,w338); //  
 nmos #(2) nmos_3_3_3_3_251_635(w340,vss,w341); //  
 pmos #(2) pmos_4_4_4_4_252_636(w340,w339,w341); //  
 nmos #(3) nmos_5_5_5_5_253_637(w34,vss,w340); //  
 pmos #(3) pmos_6_6_6_6_254_638(w34,vdd,w340); //  
 pmos #(1) pmos_1_7_7_7_255_639(w343,vdd,w342); //  
 nmos #(1) nmos_2_8_8_8_256_640(w343,vss,w342); //  
 nmos #(1) nmos_1_9_9_9_257_641(w344,vss,w343); //  
 pmos #(2) pmos_2_10_10_10_258_642(w345,vdd,w248); //  
 pmos #(2) pmos_3_11_11_11_259_643(w345,vdd,w343); //  
 nmos #(2) nmos_4_12_12_12_260_644(w345,w344,w248); //  
 nmos #(1) nmos_5_13_13_13_261_645(w338,vss,w345); //  
 pmos #(1) pmos_6_14_14_14_262_646(w338,vdd,w345); //  
 pmos #(1) pmos_1_15_15_15_263_647(w346,vdd,w248); //  
 nmos #(1) nmos_2_16_16_16_264_648(w346,vss,w248); //  
 nmos #(1) nmos_1_17_17_17_265_649(w347,vss,w346); //  
 pmos #(2) pmos_2_18_18_18_266_650(w348,vdd,w342); //  
 pmos #(2) pmos_3_19_19_19_267_651(w348,vdd,w346); //  
 nmos #(2) nmos_4_20_20_20_268_652(w348,w347,w342); //  
 nmos #(1) nmos_5_21_21_21_269_653(w341,vss,w348); //  
 pmos #(1) pmos_6_22_22_22_270_654(w341,vdd,w348); //  
 nmos #(1) nmos_1_23_23_271_655(w349,vss,w248); //  
 pmos #(2) pmos_2_24_24_272_656(w350,vdd,w342); //  
 pmos #(2) pmos_3_25_25_273_657(w350,vdd,w248); //  
 nmos #(2) nmos_4_26_26_274_658(w350,w349,w342); //  
 nmos #(1) nmos_5_27_27_275_659(w351,vss,w350); //  
 pmos #(1) pmos_6_28_28_276_660(w351,vdd,w350); //  
 pmos #(1) pmos_1_1_1_29_277_661(w353,vdd,w352); //  
 nmos #(2) nmos_2_2_2_30_278_662(w354,vss,w352); //  
 nmos #(2) nmos_3_3_3_31_279_663(w354,vss,w355); //  
 pmos #(2) pmos_4_4_4_32_280_664(w354,w353,w355); //  
 nmos #(4) nmos_5_5_5_33_281_665(w342,vss,w354); //  
 pmos #(4) pmos_6_6_6_34_282_666(w342,vdd,w354); //  
 pmos #(1) pmos_1_7_7_35_283_667(w356,vdd,w24); //  
 nmos #(1) nmos_2_8_8_36_284_668(w356,vss,w24); //  
 nmos #(1) nmos_1_9_9_37_285_669(w357,vss,w356); //  
 pmos #(2) pmos_2_10_10_38_286_670(w358,vdd,vss); //  
 pmos #(2) pmos_3_11_11_39_287_671(w358,vdd,w356); //  
 nmos #(2) nmos_4_12_12_40_288_672(w358,w357,vss); //  
 nmos #(1) nmos_5_13_13_41_289_673(w352,vss,w358); //  
 pmos #(1) pmos_6_14_14_42_290_674(w352,vdd,w358); //  
 pmos #(1) pmos_1_15_15_43_291_675(w359,vdd,vss); //  
 nmos #(1) nmos_2_16_16_44_292_676(w359,vss,vss); //  
 nmos #(1) nmos_1_17_17_45_293_677(w360,vss,w359); //  
 pmos #(2) pmos_2_18_18_46_294_678(w361,vdd,w24); //  
 pmos #(2) pmos_3_19_19_47_295_679(w361,vdd,w359); //  
 nmos #(2) nmos_4_20_20_48_296_680(w361,w360,w24); //  
 nmos #(1) nmos_5_21_21_49_297_681(w355,vss,w361); //  
 pmos #(1) pmos_6_22_22_50_298_682(w355,vdd,w361); //  
 nmos #(1) nmos_1_23_51_299_683(w362,vss,vss); //  
 pmos #(2) pmos_2_24_52_300_684(w363,vdd,w24); //  
 pmos #(2) pmos_3_25_53_301_685(w363,vdd,vss); //  
 nmos #(2) nmos_4_26_54_302_686(w363,w362,w24); //  
 nmos #(1) nmos_5_27_55_303_687(w364,vss,w363); //  
 pmos #(1) pmos_6_28_56_304_688(w364,vdd,w363); //  
 pmos #(1) pmos_1_57_305_689(w365,vdd,w364); //  
 nmos #(2) nmos_2_58_306_690(w366,vss,w364); //  
 nmos #(2) nmos_3_59_307_691(w366,vss,w351); //  
 pmos #(2) pmos_4_60_308_692(w366,w365,w351); //  
 nmos #(4) nmos_5_61_309_693(w367,vss,w366); //  
 pmos #(4) pmos_6_62_310_694(w367,vdd,w366); //  
 pmos #(1) pmos_1_1_1_1_311_695(w369,vdd,w368); //  
 nmos #(2) nmos_2_2_2_2_312_696(w370,vss,w368); //  
 nmos #(2) nmos_3_3_3_3_313_697(w370,vss,w371); //  
 pmos #(2) pmos_4_4_4_4_314_698(w370,w369,w371); //  
 nmos #(6) nmos_5_5_5_5_315_699(w33,vss,w370); //  
 pmos #(6) pmos_6_6_6_6_316_700(w33,vdd,w370); //  
 pmos #(1) pmos_1_7_7_7_317_701(w373,vdd,w372); //  
 nmos #(1) nmos_2_8_8_8_318_702(w373,vss,w372); //  
 nmos #(1) nmos_1_9_9_9_319_703(w374,vss,w373); //  
 pmos #(2) pmos_2_10_10_10_320_704(w375,vdd,w367); //  
 pmos #(2) pmos_3_11_11_11_321_705(w375,vdd,w373); //  
 nmos #(2) nmos_4_12_12_12_322_706(w375,w374,w367); //  
 nmos #(1) nmos_5_13_13_13_323_707(w368,vss,w375); //  
 pmos #(1) pmos_6_14_14_14_324_708(w368,vdd,w375); //  
 pmos #(1) pmos_1_15_15_15_325_709(w376,vdd,w367); //  
 nmos #(1) nmos_2_16_16_16_326_710(w376,vss,w367); //  
 nmos #(1) nmos_1_17_17_17_327_711(w377,vss,w376); //  
 pmos #(2) pmos_2_18_18_18_328_712(w378,vdd,w372); //  
 pmos #(2) pmos_3_19_19_19_329_713(w378,vdd,w376); //  
 nmos #(2) nmos_4_20_20_20_330_714(w378,w377,w372); //  
 nmos #(1) nmos_5_21_21_21_331_715(w371,vss,w378); //  
 pmos #(1) pmos_6_22_22_22_332_716(w371,vdd,w378); //  
 nmos #(1) nmos_1_23_23_333_717(w379,vss,w367); //  
 pmos #(2) pmos_2_24_24_334_718(w380,vdd,w372); //  
 pmos #(2) pmos_3_25_25_335_719(w380,vdd,w367); //  
 nmos #(2) nmos_4_26_26_336_720(w380,w379,w372); //  
 nmos #(1) nmos_5_27_27_337_721(w381,vss,w380); //  
 pmos #(1) pmos_6_28_28_338_722(w381,vdd,w380); //  
 pmos #(1) pmos_1_1_1_29_339_723(w383,vdd,w382); //  
 nmos #(2) nmos_2_2_2_30_340_724(w384,vss,w382); //  
 nmos #(2) nmos_3_3_3_31_341_725(w384,vss,w385); //  
 pmos #(2) pmos_4_4_4_32_342_726(w384,w383,w385); //  
 nmos #(4) nmos_5_5_5_33_343_727(w372,vss,w384); //  
 pmos #(4) pmos_6_6_6_34_344_728(w372,vdd,w384); //  
 pmos #(1) pmos_1_7_7_35_345_729(w386,vdd,w24); //  
 nmos #(1) nmos_2_8_8_36_346_730(w386,vss,w24); //  
 nmos #(1) nmos_1_9_9_37_347_731(w387,vss,w386); //  
 pmos #(2) pmos_2_10_10_38_348_732(w388,vdd,vss); //  
 pmos #(2) pmos_3_11_11_39_349_733(w388,vdd,w386); //  
 nmos #(2) nmos_4_12_12_40_350_734(w388,w387,vss); //  
 nmos #(1) nmos_5_13_13_41_351_735(w382,vss,w388); //  
 pmos #(1) pmos_6_14_14_42_352_736(w382,vdd,w388); //  
 pmos #(1) pmos_1_15_15_43_353_737(w389,vdd,vss); //  
 nmos #(1) nmos_2_16_16_44_354_738(w389,vss,vss); //  
 nmos #(1) nmos_1_17_17_45_355_739(w390,vss,w389); //  
 pmos #(2) pmos_2_18_18_46_356_740(w391,vdd,w24); //  
 pmos #(2) pmos_3_19_19_47_357_741(w391,vdd,w389); //  
 nmos #(2) nmos_4_20_20_48_358_742(w391,w390,w24); //  
 nmos #(1) nmos_5_21_21_49_359_743(w385,vss,w391); //  
 pmos #(1) pmos_6_22_22_50_360_744(w385,vdd,w391); //  
 nmos #(1) nmos_1_23_51_361_745(w392,vss,vss); //  
 pmos #(2) pmos_2_24_52_362_746(w393,vdd,w24); //  
 pmos #(2) pmos_3_25_53_363_747(w393,vdd,vss); //  
 nmos #(2) nmos_4_26_54_364_748(w393,w392,w24); //  
 nmos #(1) nmos_5_27_55_365_749(w394,vss,w393); //  
 pmos #(1) pmos_6_28_56_366_750(w394,vdd,w393); //  
 pmos #(1) pmos_1_57_367_751(w395,vdd,w394); //  
 nmos #(2) nmos_2_58_368_752(w396,vss,w394); //  
 nmos #(2) nmos_3_59_369_753(w396,vss,w381); //  
 pmos #(2) pmos_4_60_370_754(w396,w395,w381); //  
 nmos #(1) nmos_5_61_371_755(w32,vss,w396); //  
 pmos #(1) pmos_6_62_372_756(w32,vdd,w396); //  
 not #(2) NOT_1_1_757(w397,MC1);
 not #(8) NOT_2_2_758(w23,w397);
 pmos #(2) pmos_1_3_3_759(w397,vdd,MC1); //  
 nmos #(2) nmos_2_4_4_760(w397,vss,MC1); //  
 pmos #(8) pmos_1_5_5_761(w23,vdd,w397); //  
 nmos #(8) nmos_2_6_6_762(w23,vss,w397); //  
 pmos #(1) pmos_1_7_763(w399,vdd,w398); //  
 nmos #(2) nmos_2_8_764(w400,vss,w398); //  
 nmos #(2) nmos_3_9_765(w400,vss,w401); //  
 pmos #(2) pmos_4_10_766(w400,w399,w401); //  
 nmos #(3) nmos_5_11_767(w22,vss,w400); //  
 pmos #(3) pmos_6_12_768(w22,vdd,w400); //  
 pmos #(1) pmos_1_13_769(w402,vdd,MC0); //  
 nmos #(1) nmos_2_14_770(w402,vss,MC0); //  
 pmos #(1) pmos_1_1_15_771(w404,vdd,w403); //  
 nmos #(2) nmos_2_2_16_772(w405,vss,w403); //  
 nmos #(2) nmos_3_3_17_773(w405,vss,w406); //  
 pmos #(2) pmos_4_4_18_774(w405,w404,w406); //  
 nmos #(3) nmos_5_5_19_775(w21,vss,w405); //  
 pmos #(3) pmos_6_6_20_776(w21,vdd,w405); //  
 pmos #(1) pmos_1_7_21_777(w407,vdd,MC0); //  
 nmos #(1) nmos_2_8_22_778(w407,vss,MC0); //  
 nmos #(1) nmos_1_9_23_779(w408,vss,w407); //  
 pmos #(2) pmos_2_10_24_780(w409,vdd,vss); //  
 pmos #(2) pmos_3_11_25_781(w409,vdd,w407); //  
 nmos #(2) nmos_4_12_26_782(w409,w408,vss); //  
 nmos #(1) nmos_5_13_27_783(w403,vss,w409); //  
 pmos #(1) pmos_6_14_28_784(w403,vdd,w409); //  
 pmos #(1) pmos_1_15_29_785(w410,vdd,vss); //  
 nmos #(1) nmos_2_16_30_786(w410,vss,vss); //  
 nmos #(1) nmos_1_17_31_787(w411,vss,w410); //  
 pmos #(2) pmos_2_18_32_788(w412,vdd,MC0); //  
 pmos #(2) pmos_3_19_33_789(w412,vdd,w410); //  
 nmos #(2) nmos_4_20_34_790(w412,w411,MC0); //  
 nmos #(1) nmos_5_21_35_791(w406,vss,w412); //  
 pmos #(1) pmos_6_22_36_792(w406,vdd,w412); //  
 pmos #(1) pmos_1_37_793(w413,vdd,vss); //  
 nmos #(1) nmos_2_38_794(w413,vss,vss); //  
 nmos #(1) nmos_1_39_795(w414,vss,MC0); //  
 pmos #(2) pmos_2_40_796(w415,vdd,vss); //  
 pmos #(2) pmos_3_41_797(w415,vdd,MC0); //  
 nmos #(2) nmos_4_42_798(w415,w414,vss); //  
 nmos #(1) nmos_5_43_799(w416,vss,w415); //  
 pmos #(1) pmos_6_44_800(w416,vdd,w415); //  
 nmos #(1) nmos_1_45_801(w417,vss,MC1); //  
 pmos #(2) pmos_2_46_802(w419,vdd,w418); //  
 pmos #(2) pmos_3_47_803(w419,vdd,MC1); //  
 nmos #(2) nmos_4_48_804(w419,w417,w418); //  
 nmos #(1) nmos_5_49_805(w398,vss,w419); //  
 pmos #(1) pmos_6_50_806(w398,vdd,w419); //  
 nmos #(1) nmos_1_51_807(w420,vss,w402); //  
 pmos #(2) pmos_2_52_808(w421,vdd,w413); //  
 pmos #(2) pmos_3_53_809(w421,vdd,w402); //  
 nmos #(2) nmos_4_54_810(w421,w420,w413); //  
 nmos #(1) nmos_5_55_811(w418,vss,w421); //  
 pmos #(1) pmos_6_56_812(w418,vdd,w421); //  
 pmos #(1) pmos_1_57_813(w422,vdd,MC1); //  
 nmos #(1) nmos_2_58_814(w422,vss,MC1); //  
 nmos #(1) nmos_1_59_815(w423,vss,w422); //  
 pmos #(2) pmos_2_60_816(w424,vdd,w416); //  
 pmos #(2) pmos_3_61_817(w424,vdd,w422); //  
 nmos #(2) nmos_4_62_818(w424,w423,w416); //  
 nmos #(1) nmos_5_63_819(w401,vss,w424); //  
 pmos #(1) pmos_6_64_820(w401,vdd,w424); //  
 pmos #(1) pmos_1_1_1_1_1_821(w426,vdd,w425); //  
 nmos #(2) nmos_2_2_2_2_2_822(w427,vss,w425); //  
 nmos #(2) nmos_3_3_3_3_3_823(w427,vss,w428); //  
 pmos #(2) pmos_4_4_4_4_4_824(w427,w426,w428); //  
 nmos #(1) nmos_5_5_5_5_5_825(PROD5,vss,w427); //  
 pmos #(1) pmos_6_6_6_6_6_826(PROD5,vdd,w427); //  
 pmos #(1) pmos_1_7_7_7_7_827(w430,vdd,w429); //  
 nmos #(1) nmos_2_8_8_8_8_828(w430,vss,w429); //  
 nmos #(1) nmos_1_9_9_9_9_829(w431,vss,w430); //  
 pmos #(2) pmos_2_10_10_10_10_830(w433,vdd,w432); //  
 pmos #(2) pmos_3_11_11_11_11_831(w433,vdd,w430); //  
 nmos #(2) nmos_4_12_12_12_12_832(w433,w431,w432); //  
 nmos #(1) nmos_5_13_13_13_13_833(w425,vss,w433); //  
 pmos #(1) pmos_6_14_14_14_14_834(w425,vdd,w433); //  
 pmos #(1) pmos_1_15_15_15_15_835(w434,vdd,w432); //  
 nmos #(1) nmos_2_16_16_16_16_836(w434,vss,w432); //  
 nmos #(1) nmos_1_17_17_17_17_837(w435,vss,w434); //  
 pmos #(2) pmos_2_18_18_18_18_838(w436,vdd,w429); //  
 pmos #(2) pmos_3_19_19_19_19_839(w436,vdd,w434); //  
 nmos #(2) nmos_4_20_20_20_20_840(w436,w435,w429); //  
 nmos #(1) nmos_5_21_21_21_21_841(w428,vss,w436); //  
 pmos #(1) pmos_6_22_22_22_22_842(w428,vdd,w436); //  
 nmos #(1) nmos_1_23_23_23_843(w437,vss,w432); //  
 pmos #(2) pmos_2_24_24_24_844(w438,vdd,w429); //  
 pmos #(2) pmos_3_25_25_25_845(w438,vdd,w432); //  
 nmos #(2) nmos_4_26_26_26_846(w438,w437,w429); //  
 nmos #(1) nmos_5_27_27_27_847(w439,vss,w438); //  
 pmos #(1) pmos_6_28_28_28_848(w439,vdd,w438); //  
 pmos #(1) pmos_1_1_1_29_29_849(w441,vdd,w440); //  
 nmos #(2) nmos_2_2_2_30_30_850(w442,vss,w440); //  
 nmos #(2) nmos_3_3_3_31_31_851(w442,vss,w443); //  
 pmos #(2) pmos_4_4_4_32_32_852(w442,w441,w443); //  
 nmos #(4) nmos_5_5_5_33_33_853(w429,vss,w442); //  
 pmos #(4) pmos_6_6_6_34_34_854(w429,vdd,w442); //  
 pmos #(1) pmos_1_7_7_35_35_855(w444,vdd,w28); //  
 nmos #(1) nmos_2_8_8_36_36_856(w444,vss,w28); //  
 nmos #(1) nmos_1_9_9_37_37_857(w445,vss,w444); //  
 pmos #(2) pmos_2_10_10_38_38_858(w446,vdd,w33); //  
 pmos #(2) pmos_3_11_11_39_39_859(w446,vdd,w444); //  
 nmos #(2) nmos_4_12_12_40_40_860(w446,w445,w33); //  
 nmos #(1) nmos_5_13_13_41_41_861(w440,vss,w446); //  
 pmos #(1) pmos_6_14_14_42_42_862(w440,vdd,w446); //  
 pmos #(1) pmos_1_15_15_43_43_863(w447,vdd,w33); //  
 nmos #(1) nmos_2_16_16_44_44_864(w447,vss,w33); //  
 nmos #(1) nmos_1_17_17_45_45_865(w448,vss,w447); //  
 pmos #(2) pmos_2_18_18_46_46_866(w449,vdd,w28); //  
 pmos #(2) pmos_3_19_19_47_47_867(w449,vdd,w447); //  
 nmos #(2) nmos_4_20_20_48_48_868(w449,w448,w28); //  
 nmos #(1) nmos_5_21_21_49_49_869(w443,vss,w449); //  
 pmos #(1) pmos_6_22_22_50_50_870(w443,vdd,w449); //  
 nmos #(1) nmos_1_23_51_51_871(w450,vss,w33); //  
 pmos #(2) pmos_2_24_52_52_872(w451,vdd,w28); //  
 pmos #(2) pmos_3_25_53_53_873(w451,vdd,w33); //  
 nmos #(2) nmos_4_26_54_54_874(w451,w450,w28); //  
 nmos #(1) nmos_5_27_55_55_875(w452,vss,w451); //  
 pmos #(1) pmos_6_28_56_56_876(w452,vdd,w451); //  
 pmos #(1) pmos_1_57_57_877(w453,vdd,w452); //  
 nmos #(2) nmos_2_58_58_878(w454,vss,w452); //  
 nmos #(2) nmos_3_59_59_879(w454,vss,w439); //  
 pmos #(2) pmos_4_60_60_880(w454,w453,w439); //  
 nmos #(4) nmos_5_61_61_881(w455,vss,w454); //  
 pmos #(4) pmos_6_62_62_882(w455,vdd,w454); //  
 pmos #(1) pmos_1_1_1_1_63_883(w457,vdd,w456); //  
 nmos #(2) nmos_2_2_2_2_64_884(w458,vss,w456); //  
 nmos #(2) nmos_3_3_3_3_65_885(w458,vss,w459); //  
 pmos #(2) pmos_4_4_4_4_66_886(w458,w457,w459); //  
 nmos #(1) nmos_5_5_5_5_67_887(PROD2,vss,w458); //  
 pmos #(1) pmos_6_6_6_6_68_888(PROD2,vdd,w458); //  
 pmos #(1) pmos_1_7_7_7_69_889(w461,vdd,w460); //  
 nmos #(1) nmos_2_8_8_8_70_890(w461,vss,w460); //  
 nmos #(1) nmos_1_9_9_9_71_891(w462,vss,w461); //  
 pmos #(2) pmos_2_10_10_10_72_892(w463,vdd,w20); //  
 pmos #(2) pmos_3_11_11_11_73_893(w463,vdd,w461); //  
 nmos #(2) nmos_4_12_12_12_74_894(w463,w462,w20); //  
 nmos #(1) nmos_5_13_13_13_75_895(w456,vss,w463); //  
 pmos #(1) pmos_6_14_14_14_76_896(w456,vdd,w463); //  
 pmos #(1) pmos_1_15_15_15_77_897(w464,vdd,w20); //  
 nmos #(1) nmos_2_16_16_16_78_898(w464,vss,w20); //  
 nmos #(1) nmos_1_17_17_17_79_899(w465,vss,w464); //  
 pmos #(2) pmos_2_18_18_18_80_900(w466,vdd,w460); //  
 pmos #(2) pmos_3_19_19_19_81_901(w466,vdd,w464); //  
 nmos #(2) nmos_4_20_20_20_82_902(w466,w465,w460); //  
 nmos #(1) nmos_5_21_21_21_83_903(w459,vss,w466); //  
 pmos #(1) pmos_6_22_22_22_84_904(w459,vdd,w466); //  
 nmos #(1) nmos_1_23_23_85_905(w467,vss,w20); //  
 pmos #(2) pmos_2_24_24_86_906(w468,vdd,w460); //  
 pmos #(2) pmos_3_25_25_87_907(w468,vdd,w20); //  
 nmos #(2) nmos_4_26_26_88_908(w468,w467,w460); //  
 nmos #(1) nmos_5_27_27_89_909(w469,vss,w468); //  
 pmos #(1) pmos_6_28_28_90_910(w469,vdd,w468); //  
 pmos #(1) pmos_1_1_1_29_91_911(w471,vdd,w470); //  
 nmos #(2) nmos_2_2_2_30_92_912(w472,vss,w470); //  
 nmos #(2) nmos_3_3_3_31_93_913(w472,vss,w473); //  
 pmos #(2) pmos_4_4_4_32_94_914(w472,w471,w473); //  
 nmos #(4) nmos_5_5_5_33_95_915(w460,vss,w472); //  
 pmos #(4) pmos_6_6_6_34_96_916(w460,vdd,w472); //  
 pmos #(1) pmos_1_7_7_35_97_917(w474,vdd,w30); //  
 nmos #(1) nmos_2_8_8_36_98_918(w474,vss,w30); //  
 nmos #(1) nmos_1_9_9_37_99_919(w475,vss,w474); //  
 pmos #(2) pmos_2_10_10_38_100_920(w476,vdd,w36); //  
 pmos #(2) pmos_3_11_11_39_101_921(w476,vdd,w474); //  
 nmos #(2) nmos_4_12_12_40_102_922(w476,w475,w36); //  
 nmos #(1) nmos_5_13_13_41_103_923(w470,vss,w476); //  
 pmos #(1) pmos_6_14_14_42_104_924(w470,vdd,w476); //  
 pmos #(1) pmos_1_15_15_43_105_925(w477,vdd,w36); //  
 nmos #(1) nmos_2_16_16_44_106_926(w477,vss,w36); //  
 nmos #(1) nmos_1_17_17_45_107_927(w478,vss,w477); //  
 pmos #(2) pmos_2_18_18_46_108_928(w479,vdd,w30); //  
 pmos #(2) pmos_3_19_19_47_109_929(w479,vdd,w477); //  
 nmos #(2) nmos_4_20_20_48_110_930(w479,w478,w30); //  
 nmos #(1) nmos_5_21_21_49_111_931(w473,vss,w479); //  
 pmos #(1) pmos_6_22_22_50_112_932(w473,vdd,w479); //  
 nmos #(1) nmos_1_23_51_113_933(w480,vss,w36); //  
 pmos #(2) pmos_2_24_52_114_934(w481,vdd,w30); //  
 pmos #(2) pmos_3_25_53_115_935(w481,vdd,w36); //  
 nmos #(2) nmos_4_26_54_116_936(w481,w480,w30); //  
 nmos #(1) nmos_5_27_55_117_937(w482,vss,w481); //  
 pmos #(1) pmos_6_28_56_118_938(w482,vdd,w481); //  
 pmos #(1) pmos_1_57_119_939(w483,vdd,w482); //  
 nmos #(2) nmos_2_58_120_940(w484,vss,w482); //  
 nmos #(2) nmos_3_59_121_941(w484,vss,w469); //  
 pmos #(2) pmos_4_60_122_942(w484,w483,w469); //  
 nmos #(4) nmos_5_61_123_943(w485,vss,w484); //  
 pmos #(4) pmos_6_62_124_944(w485,vdd,w484); //  
 pmos #(1) pmos_1_1_1_1_125_945(w487,vdd,w486); //  
 nmos #(2) nmos_2_2_2_2_126_946(w488,vss,w486); //  
 nmos #(2) nmos_3_3_3_3_127_947(w488,vss,w489); //  
 pmos #(2) pmos_4_4_4_4_128_948(w488,w487,w489); //  
 nmos #(1) nmos_5_5_5_5_129_949(PROD3,vss,w488); //  
 pmos #(1) pmos_6_6_6_6_130_950(PROD3,vdd,w488); //  
 pmos #(1) pmos_1_7_7_7_131_951(w491,vdd,w490); //  
 nmos #(1) nmos_2_8_8_8_132_952(w491,vss,w490); //  
 nmos #(1) nmos_1_9_9_9_133_953(w492,vss,w491); //  
 pmos #(2) pmos_2_10_10_10_134_954(w493,vdd,w485); //  
 pmos #(2) pmos_3_11_11_11_135_955(w493,vdd,w491); //  
 nmos #(2) nmos_4_12_12_12_136_956(w493,w492,w485); //  
 nmos #(1) nmos_5_13_13_13_137_957(w486,vss,w493); //  
 pmos #(1) pmos_6_14_14_14_138_958(w486,vdd,w493); //  
 pmos #(1) pmos_1_15_15_15_139_959(w494,vdd,w485); //  
 nmos #(1) nmos_2_16_16_16_140_960(w494,vss,w485); //  
 nmos #(1) nmos_1_17_17_17_141_961(w495,vss,w494); //  
 pmos #(2) pmos_2_18_18_18_142_962(w496,vdd,w490); //  
 pmos #(2) pmos_3_19_19_19_143_963(w496,vdd,w494); //  
 nmos #(2) nmos_4_20_20_20_144_964(w496,w495,w490); //  
 nmos #(1) nmos_5_21_21_21_145_965(w489,vss,w496); //  
 pmos #(1) pmos_6_22_22_22_146_966(w489,vdd,w496); //  
 nmos #(1) nmos_1_23_23_147_967(w497,vss,w485); //  
 pmos #(2) pmos_2_24_24_148_968(w498,vdd,w490); //  
 pmos #(2) pmos_3_25_25_149_969(w498,vdd,w485); //  
 nmos #(2) nmos_4_26_26_150_970(w498,w497,w490); //  
 nmos #(1) nmos_5_27_27_151_971(w499,vss,w498); //  
 pmos #(1) pmos_6_28_28_152_972(w499,vdd,w498); //  
 pmos #(1) pmos_1_1_1_29_153_973(w501,vdd,w500); //  
 nmos #(2) nmos_2_2_2_30_154_974(w502,vss,w500); //  
 nmos #(2) nmos_3_3_3_31_155_975(w502,vss,w503); //  
 pmos #(2) pmos_4_4_4_32_156_976(w502,w501,w503); //  
 nmos #(4) nmos_5_5_5_33_157_977(w490,vss,w502); //  
 pmos #(4) pmos_6_6_6_34_158_978(w490,vdd,w502); //  
 pmos #(1) pmos_1_7_7_35_159_979(w504,vdd,w29); //  
 nmos #(1) nmos_2_8_8_36_160_980(w504,vss,w29); //  
 nmos #(1) nmos_1_9_9_37_161_981(w505,vss,w504); //  
 pmos #(2) pmos_2_10_10_38_162_982(w506,vdd,w35); //  
 pmos #(2) pmos_3_11_11_39_163_983(w506,vdd,w504); //  
 nmos #(2) nmos_4_12_12_40_164_984(w506,w505,w35); //  
 nmos #(1) nmos_5_13_13_41_165_985(w500,vss,w506); //  
 pmos #(1) pmos_6_14_14_42_166_986(w500,vdd,w506); //  
 pmos #(1) pmos_1_15_15_43_167_987(w507,vdd,w35); //  
 nmos #(1) nmos_2_16_16_44_168_988(w507,vss,w35); //  
 nmos #(1) nmos_1_17_17_45_169_989(w508,vss,w507); //  
 pmos #(2) pmos_2_18_18_46_170_990(w509,vdd,w29); //  
 pmos #(2) pmos_3_19_19_47_171_991(w509,vdd,w507); //  
 nmos #(2) nmos_4_20_20_48_172_992(w509,w508,w29); //  
 nmos #(1) nmos_5_21_21_49_173_993(w503,vss,w509); //  
 pmos #(1) pmos_6_22_22_50_174_994(w503,vdd,w509); //  
 nmos #(1) nmos_1_23_51_175_995(w510,vss,w35); //  
 pmos #(2) pmos_2_24_52_176_996(w511,vdd,w29); //  
 pmos #(2) pmos_3_25_53_177_997(w511,vdd,w35); //  
 nmos #(2) nmos_4_26_54_178_998(w511,w510,w29); //  
 nmos #(1) nmos_5_27_55_179_999(w512,vss,w511); //  
 pmos #(1) pmos_6_28_56_180_1000(w512,vdd,w511); //  
 pmos #(1) pmos_1_57_181_1001(w513,vdd,w512); //  
 nmos #(2) nmos_2_58_182_1002(w514,vss,w512); //  
 nmos #(2) nmos_3_59_183_1003(w514,vss,w499); //  
 pmos #(2) pmos_4_60_184_1004(w514,w513,w499); //  
 nmos #(4) nmos_5_61_185_1005(w515,vss,w514); //  
 pmos #(4) pmos_6_62_186_1006(w515,vdd,w514); //  
 pmos #(1) pmos_1_1_1_1_187_1007(w517,vdd,w516); //  
 nmos #(2) nmos_2_2_2_2_188_1008(w518,vss,w516); //  
 nmos #(2) nmos_3_3_3_3_189_1009(w518,vss,w519); //  
 pmos #(2) pmos_4_4_4_4_190_1010(w518,w517,w519); //  
 nmos #(1) nmos_5_5_5_5_191_1011(PROD4,vss,w518); //  
 pmos #(1) pmos_6_6_6_6_192_1012(PROD4,vdd,w518); //  
 pmos #(1) pmos_1_7_7_7_193_1013(w521,vdd,w520); //  
 nmos #(1) nmos_2_8_8_8_194_1014(w521,vss,w520); //  
 nmos #(1) nmos_1_9_9_9_195_1015(w522,vss,w521); //  
 pmos #(2) pmos_2_10_10_10_196_1016(w523,vdd,w515); //  
 pmos #(2) pmos_3_11_11_11_197_1017(w523,vdd,w521); //  
 nmos #(2) nmos_4_12_12_12_198_1018(w523,w522,w515); //  
 nmos #(1) nmos_5_13_13_13_199_1019(w516,vss,w523); //  
 pmos #(1) pmos_6_14_14_14_200_1020(w516,vdd,w523); //  
 pmos #(1) pmos_1_15_15_15_201_1021(w524,vdd,w515); //  
 nmos #(1) nmos_2_16_16_16_202_1022(w524,vss,w515); //  
 nmos #(1) nmos_1_17_17_17_203_1023(w525,vss,w524); //  
 pmos #(2) pmos_2_18_18_18_204_1024(w526,vdd,w520); //  
 pmos #(2) pmos_3_19_19_19_205_1025(w526,vdd,w524); //  
 nmos #(2) nmos_4_20_20_20_206_1026(w526,w525,w520); //  
 nmos #(1) nmos_5_21_21_21_207_1027(w519,vss,w526); //  
 pmos #(1) pmos_6_22_22_22_208_1028(w519,vdd,w526); //  
 nmos #(1) nmos_1_23_23_209_1029(w527,vss,w515); //  
 pmos #(2) pmos_2_24_24_210_1030(w528,vdd,w520); //  
 pmos #(2) pmos_3_25_25_211_1031(w528,vdd,w515); //  
 nmos #(2) nmos_4_26_26_212_1032(w528,w527,w520); //  
 nmos #(1) nmos_5_27_27_213_1033(w529,vss,w528); //  
 pmos #(1) pmos_6_28_28_214_1034(w529,vdd,w528); //  
 pmos #(1) pmos_1_1_1_29_215_1035(w531,vdd,w530); //  
 nmos #(2) nmos_2_2_2_30_216_1036(w532,vss,w530); //  
 nmos #(2) nmos_3_3_3_31_217_1037(w532,vss,w533); //  
 pmos #(2) pmos_4_4_4_32_218_1038(w532,w531,w533); //  
 nmos #(4) nmos_5_5_5_33_219_1039(w520,vss,w532); //  
 pmos #(4) pmos_6_6_6_34_220_1040(w520,vdd,w532); //  
 pmos #(1) pmos_1_7_7_35_221_1041(w534,vdd,w31); //  
 nmos #(1) nmos_2_8_8_36_222_1042(w534,vss,w31); //  
 nmos #(1) nmos_1_9_9_37_223_1043(w535,vss,w534); //  
 pmos #(2) pmos_2_10_10_38_224_1044(w536,vdd,w34); //  
 pmos #(2) pmos_3_11_11_39_225_1045(w536,vdd,w534); //  
 nmos #(2) nmos_4_12_12_40_226_1046(w536,w535,w34); //  
 nmos #(1) nmos_5_13_13_41_227_1047(w530,vss,w536); //  
 pmos #(1) pmos_6_14_14_42_228_1048(w530,vdd,w536); //  
 pmos #(1) pmos_1_15_15_43_229_1049(w537,vdd,w34); //  
 nmos #(1) nmos_2_16_16_44_230_1050(w537,vss,w34); //  
 nmos #(1) nmos_1_17_17_45_231_1051(w538,vss,w537); //  
 pmos #(2) pmos_2_18_18_46_232_1052(w539,vdd,w31); //  
 pmos #(2) pmos_3_19_19_47_233_1053(w539,vdd,w537); //  
 nmos #(2) nmos_4_20_20_48_234_1054(w539,w538,w31); //  
 nmos #(1) nmos_5_21_21_49_235_1055(w533,vss,w539); //  
 pmos #(1) pmos_6_22_22_50_236_1056(w533,vdd,w539); //  
 nmos #(1) nmos_1_23_51_237_1057(w540,vss,w34); //  
 pmos #(2) pmos_2_24_52_238_1058(w541,vdd,w31); //  
 pmos #(2) pmos_3_25_53_239_1059(w541,vdd,w34); //  
 nmos #(2) nmos_4_26_54_240_1060(w541,w540,w31); //  
 nmos #(1) nmos_5_27_55_241_1061(w542,vss,w541); //  
 pmos #(1) pmos_6_28_56_242_1062(w542,vdd,w541); //  
 pmos #(1) pmos_1_57_243_1063(w543,vdd,w542); //  
 nmos #(2) nmos_2_58_244_1064(w544,vss,w542); //  
 nmos #(2) nmos_3_59_245_1065(w544,vss,w529); //  
 pmos #(2) pmos_4_60_246_1066(w544,w543,w529); //  
 nmos #(4) nmos_5_61_247_1067(w432,vss,w544); //  
 pmos #(4) pmos_6_62_248_1068(w432,vdd,w544); //  
 pmos #(1) pmos_1_1_1_1_249_1069(w546,vdd,w545); //  
 nmos #(2) nmos_2_2_2_2_250_1070(w547,vss,w545); //  
 nmos #(2) nmos_3_3_3_3_251_1071(w547,vss,w548); //  
 pmos #(2) pmos_4_4_4_4_252_1072(w547,w546,w548); //  
 nmos #(1) nmos_5_5_5_5_253_1073(PROD6,vss,w547); //  
 pmos #(1) pmos_6_6_6_6_254_1074(PROD6,vdd,w547); //  
 pmos #(1) pmos_1_7_7_7_255_1075(w550,vdd,w549); //  
 nmos #(1) nmos_2_8_8_8_256_1076(w550,vss,w549); //  
 nmos #(1) nmos_1_9_9_9_257_1077(w551,vss,w550); //  
 pmos #(2) pmos_2_10_10_10_258_1078(w552,vdd,w455); //  
 pmos #(2) pmos_3_11_11_11_259_1079(w552,vdd,w550); //  
 nmos #(2) nmos_4_12_12_12_260_1080(w552,w551,w455); //  
 nmos #(1) nmos_5_13_13_13_261_1081(w545,vss,w552); //  
 pmos #(1) pmos_6_14_14_14_262_1082(w545,vdd,w552); //  
 pmos #(1) pmos_1_15_15_15_263_1083(w553,vdd,w455); //  
 nmos #(1) nmos_2_16_16_16_264_1084(w553,vss,w455); //  
 nmos #(1) nmos_1_17_17_17_265_1085(w554,vss,w553); //  
 pmos #(2) pmos_2_18_18_18_266_1086(w555,vdd,w549); //  
 pmos #(2) pmos_3_19_19_19_267_1087(w555,vdd,w553); //  
 nmos #(2) nmos_4_20_20_20_268_1088(w555,w554,w549); //  
 nmos #(1) nmos_5_21_21_21_269_1089(w548,vss,w555); //  
 pmos #(1) pmos_6_22_22_22_270_1090(w548,vdd,w555); //  
 nmos #(1) nmos_1_23_23_271_1091(w556,vss,w455); //  
 pmos #(2) pmos_2_24_24_272_1092(w557,vdd,w549); //  
 pmos #(2) pmos_3_25_25_273_1093(w557,vdd,w455); //  
 nmos #(2) nmos_4_26_26_274_1094(w557,w556,w549); //  
 nmos #(1) nmos_5_27_27_275_1095(w558,vss,w557); //  
 pmos #(1) pmos_6_28_28_276_1096(w558,vdd,w557); //  
 pmos #(1) pmos_1_1_1_29_277_1097(w560,vdd,w559); //  
 nmos #(2) nmos_2_2_2_30_278_1098(w561,vss,w559); //  
 nmos #(2) nmos_3_3_3_31_279_1099(w561,vss,w562); //  
 pmos #(2) pmos_4_4_4_32_280_1100(w561,w560,w562); //  
 nmos #(4) nmos_5_5_5_33_281_1101(w549,vss,w561); //  
 pmos #(4) pmos_6_6_6_34_282_1102(w549,vdd,w561); //  
 pmos #(1) pmos_1_7_7_35_283_1103(w563,vdd,w28); //  
 nmos #(1) nmos_2_8_8_36_284_1104(w563,vss,w28); //  
 nmos #(1) nmos_1_9_9_37_285_1105(w564,vss,w563); //  
 pmos #(2) pmos_2_10_10_38_286_1106(w565,vdd,w33); //  
 pmos #(2) pmos_3_11_11_39_287_1107(w565,vdd,w563); //  
 nmos #(2) nmos_4_12_12_40_288_1108(w565,w564,w33); //  
 nmos #(1) nmos_5_13_13_41_289_1109(w559,vss,w565); //  
 pmos #(1) pmos_6_14_14_42_290_1110(w559,vdd,w565); //  
 pmos #(1) pmos_1_15_15_43_291_1111(w566,vdd,w33); //  
 nmos #(1) nmos_2_16_16_44_292_1112(w566,vss,w33); //  
 nmos #(1) nmos_1_17_17_45_293_1113(w567,vss,w566); //  
 pmos #(2) pmos_2_18_18_46_294_1114(w568,vdd,w28); //  
 pmos #(2) pmos_3_19_19_47_295_1115(w568,vdd,w566); //  
 nmos #(2) nmos_4_20_20_48_296_1116(w568,w567,w28); //  
 nmos #(1) nmos_5_21_21_49_297_1117(w562,vss,w568); //  
 pmos #(1) pmos_6_22_22_50_298_1118(w562,vdd,w568); //  
 nmos #(1) nmos_1_23_51_299_1119(w569,vss,w33); //  
 pmos #(2) pmos_2_24_52_300_1120(w570,vdd,w28); //  
 pmos #(2) pmos_3_25_53_301_1121(w570,vdd,w33); //  
 nmos #(2) nmos_4_26_54_302_1122(w570,w569,w28); //  
 nmos #(1) nmos_5_27_55_303_1123(w571,vss,w570); //  
 pmos #(1) pmos_6_28_56_304_1124(w571,vdd,w570); //  
 pmos #(1) pmos_1_57_305_1125(w572,vdd,w571); //  
 nmos #(2) nmos_2_58_306_1126(w573,vss,w571); //  
 nmos #(2) nmos_3_59_307_1127(w573,vss,w558); //  
 pmos #(2) pmos_4_60_308_1128(w573,w572,w558); //  
 nmos #(4) nmos_5_61_309_1129(w574,vss,w573); //  
 pmos #(4) pmos_6_62_310_1130(w574,vdd,w573); //  
 pmos #(1) pmos_1_1_1_1_311_1131(w576,vdd,w575); //  
 nmos #(2) nmos_2_2_2_2_312_1132(w577,vss,w575); //  
 nmos #(2) nmos_3_3_3_3_313_1133(w577,vss,w578); //  
 pmos #(2) pmos_4_4_4_4_314_1134(w577,w576,w578); //  
 nmos #(1) nmos_5_5_5_5_315_1135(PROD7,vss,w577); //  
 pmos #(1) pmos_6_6_6_6_316_1136(PROD7,vdd,w577); //  
 pmos #(1) pmos_1_7_7_7_317_1137(w580,vdd,w579); //  
 nmos #(1) nmos_2_8_8_8_318_1138(w580,vss,w579); //  
 nmos #(1) nmos_1_9_9_9_319_1139(w581,vss,w580); //  
 pmos #(2) pmos_2_10_10_10_320_1140(w582,vdd,w574); //  
 pmos #(2) pmos_3_11_11_11_321_1141(w582,vdd,w580); //  
 nmos #(2) nmos_4_12_12_12_322_1142(w582,w581,w574); //  
 nmos #(1) nmos_5_13_13_13_323_1143(w575,vss,w582); //  
 pmos #(1) pmos_6_14_14_14_324_1144(w575,vdd,w582); //  
 pmos #(1) pmos_1_15_15_15_325_1145(w583,vdd,w574); //  
 nmos #(1) nmos_2_16_16_16_326_1146(w583,vss,w574); //  
 nmos #(1) nmos_1_17_17_17_327_1147(w584,vss,w583); //  
 pmos #(2) pmos_2_18_18_18_328_1148(w585,vdd,w579); //  
 pmos #(2) pmos_3_19_19_19_329_1149(w585,vdd,w583); //  
 nmos #(2) nmos_4_20_20_20_330_1150(w585,w584,w579); //  
 nmos #(1) nmos_5_21_21_21_331_1151(w578,vss,w585); //  
 pmos #(1) pmos_6_22_22_22_332_1152(w578,vdd,w585); //  
 nmos #(1) nmos_1_23_23_333_1153(w586,vss,w574); //  
 pmos #(2) pmos_2_24_24_334_1154(w587,vdd,w579); //  
 pmos #(2) pmos_3_25_25_335_1155(w587,vdd,w574); //  
 nmos #(2) nmos_4_26_26_336_1156(w587,w586,w579); //  
 nmos #(1) nmos_5_27_27_337_1157(w588,vss,w587); //  
 pmos #(1) pmos_6_28_28_338_1158(w588,vdd,w587); //  
 pmos #(1) pmos_1_1_1_29_339_1159(w590,vdd,w589); //  
 nmos #(2) nmos_2_2_2_30_340_1160(w591,vss,w589); //  
 nmos #(2) nmos_3_3_3_31_341_1161(w591,vss,w592); //  
 pmos #(2) pmos_4_4_4_32_342_1162(w591,w590,w592); //  
 nmos #(4) nmos_5_5_5_33_343_1163(w579,vss,w591); //  
 pmos #(4) pmos_6_6_6_34_344_1164(w579,vdd,w591); //  
 pmos #(1) pmos_1_7_7_35_345_1165(w593,vdd,w28); //  
 nmos #(1) nmos_2_8_8_36_346_1166(w593,vss,w28); //  
 nmos #(1) nmos_1_9_9_37_347_1167(w594,vss,w593); //  
 pmos #(2) pmos_2_10_10_38_348_1168(w595,vdd,w33); //  
 pmos #(2) pmos_3_11_11_39_349_1169(w595,vdd,w593); //  
 nmos #(2) nmos_4_12_12_40_350_1170(w595,w594,w33); //  
 nmos #(1) nmos_5_13_13_41_351_1171(w589,vss,w595); //  
 pmos #(1) pmos_6_14_14_42_352_1172(w589,vdd,w595); //  
 pmos #(1) pmos_1_15_15_43_353_1173(w596,vdd,w33); //  
 nmos #(1) nmos_2_16_16_44_354_1174(w596,vss,w33); //  
 nmos #(1) nmos_1_17_17_45_355_1175(w597,vss,w596); //  
 pmos #(2) pmos_2_18_18_46_356_1176(w598,vdd,w28); //  
 pmos #(2) pmos_3_19_19_47_357_1177(w598,vdd,w596); //  
 nmos #(2) nmos_4_20_20_48_358_1178(w598,w597,w28); //  
 nmos #(1) nmos_5_21_21_49_359_1179(w592,vss,w598); //  
 pmos #(1) pmos_6_22_22_50_360_1180(w592,vdd,w598); //  
 nmos #(1) nmos_1_23_51_361_1181(w599,vss,w33); //  
 pmos #(2) pmos_2_24_52_362_1182(w600,vdd,w28); //  
 pmos #(2) pmos_3_25_53_363_1183(w600,vdd,w33); //  
 nmos #(2) nmos_4_26_54_364_1184(w600,w599,w28); //  
 nmos #(1) nmos_5_27_55_365_1185(w601,vss,w600); //  
 pmos #(1) pmos_6_28_56_366_1186(w601,vdd,w600); //  
 pmos #(1) pmos_1_57_367_1187(w602,vdd,w601); //  
 nmos #(2) nmos_2_58_368_1188(w603,vss,w601); //  
 nmos #(2) nmos_3_59_369_1189(w603,vss,w588); //  
 pmos #(2) pmos_4_60_370_1190(w603,w602,w588); //  
 nmos #(1) nmos_5_61_371_1191(w37,vss,w603); //  
 pmos #(1) pmos_6_62_372_1192(w37,vdd,w603); //  
endmodule

// Simulation parameters in Verilog Format
always
#200 MC3=~MC3;
#400 MC2=~MC2;
#800 MC1=~MC1;
#1600 MC0=~MC0;
#3200 MP3=~MP3;
#6400 MP2=~MP2;
#12800 MP1=~MP1;
#25600 MP0=~MP0;

// Simulation parameters
// MC3 CLK 1 1
// MC2 CLK 2 2
// MC1 CLK 4 4
// MC0 CLK 8 8
// MP3 CLK 16 16
// MP2 CLK 32 32
// MP1 CLK 64 64
// MP0 CLK 128 128
